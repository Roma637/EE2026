`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12.04.2025 11:02:29
// Design Name: 
// Module Name: draw_menu
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module shiftColor(
    input  [15:0] color,
    output [15:0] outputColor
);
    assign outputColor = {
        (color[15:11] >> 1), 
        (color[10:5]  >> 1), 
        (color[4:0]   >> 1)
    };
endmodule

module draw_menu(
    input clk,
    input [7:0] x,
    input [6:0] y,
    input [1:0] item_1_id,
    input [1:0] item_2_id,
    input [1:0] item_3_id,
    input [15:0] sw,
    output reg [15:0] oled_data,
    input [11:0] inventory,
    input [2:0] orders_done
);


parameter FRAME_WIDTH  = 96;
parameter FRAME_HEIGHT = 64;


wire [7:0] rot_x = FRAME_WIDTH  - 1 - x;
wire [6:0] rot_y = FRAME_HEIGHT - 1 - y;

wire [11:0] holding_ingredient_id;
assign holding_ingredient_id = inventory;


reg [15:0] chicken_rice  [0:31][0:31];
reg [15:0] onion_soup    [0:31][0:31];
reg [15:0] tomato_soup   [0:31][0:31];
reg [15:0] tomato_rice   [0:31][0:31];
reg [15:0] chicken_rice_dim  [0:31][0:31];
reg [15:0] onion_soup_dim    [0:31][0:31];
reg [15:0] tomato_soup_dim   [0:31][0:31];
reg [15:0] tomato_rice_dim   [0:31][0:31];
reg [15:0] tick_overlay   [0:31][0:31];
reg [15:0] ingredient_text [0:16][0:79];

reg [15:0] cross                  [0:14][0:14];
reg [15:0] rice_raw               [0:14][0:14];
reg [15:0] rice_boiled            [0:14][0:14];
reg [15:0] rice_chopped           [0:14][0:14];
reg [15:0] rice_boiled_chopped    [0:14][0:14];
reg [15:0] tomato_raw             [0:14][0:14];
reg [15:0] tomato_boiled          [0:14][0:14];
reg [15:0] tomato_chopped         [0:14][0:14];
reg [15:0] tomato_boiled_chopped  [0:14][0:14];
reg [15:0] chicken_raw            [0:14][0:14];
reg [15:0] chicken_boiled         [0:14][0:14];
reg [15:0] chicken_chopped        [0:14][0:14];
reg [15:0] chicken_boiled_chopped [0:14][0:14];
reg [15:0] onion_raw              [0:14][0:14];
reg [15:0] onion_boiled           [0:14][0:14];
reg [15:0] onion_chopped          [0:14][0:14];
reg [15:0] onion_boiled_chopped   [0:14][0:14];




reg [7:0] item_1_x_offset = 0;
reg [6:0] item_1_y_offset = 0;

reg [7:0] item_2_x_offset = 32;
reg [6:0] item_2_y_offset = 0;

reg [7:0] item_3_x_offset = 64;
reg [6:0] item_3_y_offset = 0;


reg [7:0] ingredient_text_x_offset = 0;
reg [6:0] ingredient_text_y_offset = 47;


reg [7:0] holding_ingredient_x_offset = 80;
reg [6:0] holding_ingredient_y_offset = 49;


reg [7:0] item_1_ingredient_1_x_offset = 1;
reg [6:0] item_1_ingredient_1_y_offset = 32;

reg [7:0] item_1_ingredient_2_x_offset = 16;
reg [6:0] item_1_ingredient_2_y_offset = 32;

reg [7:0] item_2_ingredient_1_x_offset = 33;
reg [6:0] item_2_ingredient_1_y_offset = 32;

reg [7:0] item_2_ingredient_2_x_offset = 49;
reg [6:0] item_2_ingredient_2_y_offset = 32;

reg [7:0] item_3_ingredient_1_x_offset = 65;
reg [6:0] item_3_ingredient_1_y_offset = 32;

reg [7:0] item_3_ingredient_2_x_offset = 80;
reg [6:0] item_3_ingredient_2_y_offset = 32;

//======================================================================
// Bunch of sprites
initial begin
        cross[0][0] = 16'b11111_101001_10100;
        cross[0][1] = 16'b11111_101001_10100;
        cross[0][2] = 16'b11111_101001_10100;
        cross[0][3] = 16'b11111_101001_10100;
        cross[0][4] = 16'b11111_101001_10100;
        cross[0][5] = 16'b11111_101001_10100;
        cross[0][6] = 16'b11111_101001_10100;
        cross[0][7] = 16'b11111_101001_10100;
        cross[0][8] = 16'b11111_101001_10100;
        cross[0][9] = 16'b11111_101001_10100;
        cross[0][10] = 16'b11111_101001_10100;
        cross[0][11] = 16'b11111_101001_10100;
        cross[0][12] = 16'b11111_101001_10100;
        cross[0][13] = 16'b11111_101001_10100;
        cross[0][14] = 16'b11111_101001_10100;
        cross[1][0] = 16'b11111_101001_10100;
        cross[1][1] = 16'b00000_000000_00000;
        cross[1][2] = 16'b00000_000000_00000;
        cross[1][3] = 16'b00000_000000_00000;
        cross[1][4] = 16'b00000_000000_00000;
        cross[1][5] = 16'b00000_000000_00000;
        cross[1][6] = 16'b00000_000000_00000;
        cross[1][7] = 16'b00000_000000_00000;
        cross[1][8] = 16'b00000_000000_00000;
        cross[1][9] = 16'b00000_000000_00000;
        cross[1][10] = 16'b00000_000000_00000;
        cross[1][11] = 16'b00000_000000_00000;
        cross[1][12] = 16'b00000_000000_00000;
        cross[1][13] = 16'b00000_000000_00000;
        cross[1][14] = 16'b11111_101001_10100;
        cross[2][0] = 16'b11111_101001_10100;
        cross[2][1] = 16'b00000_000000_00000;
        cross[2][2] = 16'b11111_101001_10100;
        cross[2][3] = 16'b11111_101001_10100;
        cross[2][4] = 16'b00000_000000_00000;
        cross[2][5] = 16'b00000_000000_00000;
        cross[2][6] = 16'b00000_000000_00000;
        cross[2][7] = 16'b00000_000000_00000;
        cross[2][8] = 16'b00000_000000_00000;
        cross[2][9] = 16'b00000_000000_00000;
        cross[2][10] = 16'b00000_000000_00000;
        cross[2][11] = 16'b11111_101001_10100;
        cross[2][12] = 16'b11111_101001_10100;
        cross[2][13] = 16'b00000_000000_00000;
        cross[2][14] = 16'b11111_101001_10100;
        cross[3][0] = 16'b11111_101001_10100;
        cross[3][1] = 16'b00000_000000_00000;
        cross[3][2] = 16'b11111_101001_10100;
        cross[3][3] = 16'b11111_101001_10100;
        cross[3][4] = 16'b11111_101001_10100;
        cross[3][5] = 16'b00000_000000_00000;
        cross[3][6] = 16'b00000_000000_00000;
        cross[3][7] = 16'b00000_000000_00000;
        cross[3][8] = 16'b00000_000000_00000;
        cross[3][9] = 16'b00000_000000_00000;
        cross[3][10] = 16'b11111_101001_10100;
        cross[3][11] = 16'b11111_101001_10100;
        cross[3][12] = 16'b11111_101001_10100;
        cross[3][13] = 16'b00000_000000_00000;
        cross[3][14] = 16'b11111_101001_10100;
        cross[4][0] = 16'b11111_101001_10100;
        cross[4][1] = 16'b00000_000000_00000;
        cross[4][2] = 16'b00000_000000_00000;
        cross[4][3] = 16'b11111_101001_10100;
        cross[4][4] = 16'b11111_101001_10100;
        cross[4][5] = 16'b11111_101001_10100;
        cross[4][6] = 16'b00000_000000_00000;
        cross[4][7] = 16'b00000_000000_00000;
        cross[4][8] = 16'b00000_000000_00000;
        cross[4][9] = 16'b11111_101001_10100;
        cross[4][10] = 16'b11111_101001_10100;
        cross[4][11] = 16'b11111_101001_10100;
        cross[4][12] = 16'b00000_000000_00000;
        cross[4][13] = 16'b00000_000000_00000;
        cross[4][14] = 16'b11111_101001_10100;
        cross[5][0] = 16'b11111_101001_10100;
        cross[5][1] = 16'b00000_000000_00000;
        cross[5][2] = 16'b00000_000000_00000;
        cross[5][3] = 16'b00000_000000_00000;
        cross[5][4] = 16'b11111_101001_10100;
        cross[5][5] = 16'b11111_101001_10100;
        cross[5][6] = 16'b11111_101001_10100;
        cross[5][7] = 16'b00000_000000_00000;
        cross[5][8] = 16'b11111_101001_10100;
        cross[5][9] = 16'b11111_101001_10100;
        cross[5][10] = 16'b11111_101001_10100;
        cross[5][11] = 16'b00000_000000_00000;
        cross[5][12] = 16'b00000_000000_00000;
        cross[5][13] = 16'b00000_000000_00000;
        cross[5][14] = 16'b11111_101001_10100;
        cross[6][0] = 16'b11111_101001_10100;
        cross[6][1] = 16'b00000_000000_00000;
        cross[6][2] = 16'b00000_000000_00000;
        cross[6][3] = 16'b00000_000000_00000;
        cross[6][4] = 16'b00000_000000_00000;
        cross[6][5] = 16'b11111_101001_10100;
        cross[6][6] = 16'b11111_101001_10100;
        cross[6][7] = 16'b11111_101001_10100;
        cross[6][8] = 16'b11111_101001_10100;
        cross[6][9] = 16'b11111_101001_10100;
        cross[6][10] = 16'b00000_000000_00000;
        cross[6][11] = 16'b00000_000000_00000;
        cross[6][12] = 16'b00000_000000_00000;
        cross[6][13] = 16'b00000_000000_00000;
        cross[6][14] = 16'b11111_101001_10100;
        cross[7][0] = 16'b11111_101001_10100;
        cross[7][1] = 16'b00000_000000_00000;
        cross[7][2] = 16'b00000_000000_00000;
        cross[7][3] = 16'b00000_000000_00000;
        cross[7][4] = 16'b00000_000000_00000;
        cross[7][5] = 16'b00000_000000_00000;
        cross[7][6] = 16'b11111_101001_10100;
        cross[7][7] = 16'b11111_101001_10100;
        cross[7][8] = 16'b11111_101001_10100;
        cross[7][9] = 16'b00000_000000_00000;
        cross[7][10] = 16'b00000_000000_00000;
        cross[7][11] = 16'b00000_000000_00000;
        cross[7][12] = 16'b00000_000000_00000;
        cross[7][13] = 16'b00000_000000_00000;
        cross[7][14] = 16'b11111_101001_10100;
        cross[8][0] = 16'b11111_101001_10100;
        cross[8][1] = 16'b00000_000000_00000;
        cross[8][2] = 16'b00000_000000_00000;
        cross[8][3] = 16'b00000_000000_00000;
        cross[8][4] = 16'b00000_000000_00000;
        cross[8][5] = 16'b11111_101001_10100;
        cross[8][6] = 16'b11111_101001_10100;
        cross[8][7] = 16'b11111_101001_10100;
        cross[8][8] = 16'b11111_101001_10100;
        cross[8][9] = 16'b11111_101001_10100;
        cross[8][10] = 16'b00000_000000_00000;
        cross[8][11] = 16'b00000_000000_00000;
        cross[8][12] = 16'b00000_000000_00000;
        cross[8][13] = 16'b00000_000000_00000;
        cross[8][14] = 16'b11111_101001_10100;
        cross[9][0] = 16'b11111_101001_10100;
        cross[9][1] = 16'b00000_000000_00000;
        cross[9][2] = 16'b00000_000000_00000;
        cross[9][3] = 16'b00000_000000_00000;
        cross[9][4] = 16'b11111_101001_10100;
        cross[9][5] = 16'b11111_101001_10100;
        cross[9][6] = 16'b11111_101001_10100;
        cross[9][7] = 16'b00000_000000_00000;
        cross[9][8] = 16'b11111_101001_10100;
        cross[9][9] = 16'b11111_101001_10100;
        cross[9][10] = 16'b11111_101001_10100;
        cross[9][11] = 16'b00000_000000_00000;
        cross[9][12] = 16'b00000_000000_00000;
        cross[9][13] = 16'b00000_000000_00000;
        cross[9][14] = 16'b11111_101001_10100;
        cross[10][0] = 16'b11111_101001_10100;
        cross[10][1] = 16'b00000_000000_00000;
        cross[10][2] = 16'b00000_000000_00000;
        cross[10][3] = 16'b11111_101001_10100;
        cross[10][4] = 16'b11111_101001_10100;
        cross[10][5] = 16'b11111_101001_10100;
        cross[10][6] = 16'b00000_000000_00000;
        cross[10][7] = 16'b00000_000000_00000;
        cross[10][8] = 16'b00000_000000_00000;
        cross[10][9] = 16'b11111_101001_10100;
        cross[10][10] = 16'b11111_101001_10100;
        cross[10][11] = 16'b11111_101001_10100;
        cross[10][12] = 16'b00000_000000_00000;
        cross[10][13] = 16'b00000_000000_00000;
        cross[10][14] = 16'b11111_101001_10100;
        cross[11][0] = 16'b11111_101001_10100;
        cross[11][1] = 16'b00000_000000_00000;
        cross[11][2] = 16'b11111_101001_10100;
        cross[11][3] = 16'b11111_101001_10100;
        cross[11][4] = 16'b11111_101001_10100;
        cross[11][5] = 16'b00000_000000_00000;
        cross[11][6] = 16'b00000_000000_00000;
        cross[11][7] = 16'b00000_000000_00000;
        cross[11][8] = 16'b00000_000000_00000;
        cross[11][9] = 16'b00000_000000_00000;
        cross[11][10] = 16'b11111_101001_10100;
        cross[11][11] = 16'b11111_101001_10100;
        cross[11][12] = 16'b11111_101001_10100;
        cross[11][13] = 16'b00000_000000_00000;
        cross[11][14] = 16'b11111_101001_10100;
        cross[12][0] = 16'b11111_101001_10100;
        cross[12][1] = 16'b00000_000000_00000;
        cross[12][2] = 16'b11111_101001_10100;
        cross[12][3] = 16'b11111_101001_10100;
        cross[12][4] = 16'b00000_000000_00000;
        cross[12][5] = 16'b00000_000000_00000;
        cross[12][6] = 16'b00000_000000_00000;
        cross[12][7] = 16'b00000_000000_00000;
        cross[12][8] = 16'b00000_000000_00000;
        cross[12][9] = 16'b00000_000000_00000;
        cross[12][10] = 16'b00000_000000_00000;
        cross[12][11] = 16'b11111_101001_10100;
        cross[12][12] = 16'b11111_101001_10100;
        cross[12][13] = 16'b00000_000000_00000;
        cross[12][14] = 16'b11111_101001_10100;
        cross[13][0] = 16'b11111_101001_10100;
        cross[13][1] = 16'b00000_000000_00000;
        cross[13][2] = 16'b00000_000000_00000;
        cross[13][3] = 16'b00000_000000_00000;
        cross[13][4] = 16'b00000_000000_00000;
        cross[13][5] = 16'b00000_000000_00000;
        cross[13][6] = 16'b00000_000000_00000;
        cross[13][7] = 16'b00000_000000_00000;
        cross[13][8] = 16'b00000_000000_00000;
        cross[13][9] = 16'b00000_000000_00000;
        cross[13][10] = 16'b00000_000000_00000;
        cross[13][11] = 16'b00000_000000_00000;
        cross[13][12] = 16'b00000_000000_00000;
        cross[13][13] = 16'b00000_000000_00000;
        cross[13][14] = 16'b11111_101001_10100;
        cross[14][0] = 16'b11111_101001_10100;
        cross[14][1] = 16'b11111_101001_10100;
        cross[14][2] = 16'b11111_101001_10100;
        cross[14][3] = 16'b11111_101001_10100;
        cross[14][4] = 16'b11111_101001_10100;
        cross[14][5] = 16'b11111_101001_10100;
        cross[14][6] = 16'b11111_101001_10100;
        cross[14][7] = 16'b11111_101001_10100;
        cross[14][8] = 16'b11111_101001_10100;
        cross[14][9] = 16'b11111_101001_10100;
        cross[14][10] = 16'b11111_101001_10100;
        cross[14][11] = 16'b11111_101001_10100;
        cross[14][12] = 16'b11111_101001_10100;
        cross[14][13] = 16'b11111_101001_10100;
        cross[14][14] = 16'b11111_101001_10100;


        chicken_rice[0][0] = 16'b10111_110111_11111;
        chicken_rice[0][1] = 16'b10111_110111_11111;
        chicken_rice[0][2] = 16'b10111_110111_11111;
        chicken_rice[0][3] = 16'b10111_110111_11111;
        chicken_rice[0][4] = 16'b10111_110111_11111;
        chicken_rice[0][5] = 16'b10111_110111_11111;
        chicken_rice[0][6] = 16'b10111_110111_11111;
        chicken_rice[0][7] = 16'b10111_110111_11111;
        chicken_rice[0][8] = 16'b10111_110111_11111;
        chicken_rice[0][9] = 16'b10111_110111_11111;
        chicken_rice[0][10] = 16'b10111_110111_11111;
        chicken_rice[0][11] = 16'b10111_110111_11111;
        chicken_rice[0][12] = 16'b10111_110111_11111;
        chicken_rice[0][13] = 16'b10111_110111_11111;
        chicken_rice[0][14] = 16'b10111_110111_11111;
        chicken_rice[0][15] = 16'b10111_110111_11111;
        chicken_rice[0][16] = 16'b10111_110111_11111;
        chicken_rice[0][17] = 16'b10111_110111_11111;
        chicken_rice[0][18] = 16'b10111_110111_11111;
        chicken_rice[0][19] = 16'b10111_110111_11111;
        chicken_rice[0][20] = 16'b10111_110111_11111;
        chicken_rice[0][21] = 16'b10111_110111_11111;
        chicken_rice[0][22] = 16'b10111_110111_11111;
        chicken_rice[0][23] = 16'b10111_110111_11111;
        chicken_rice[0][24] = 16'b10111_110111_11111;
        chicken_rice[0][25] = 16'b10111_110111_11111;
        chicken_rice[0][26] = 16'b10111_110111_11111;
        chicken_rice[0][27] = 16'b10111_110111_11111;
        chicken_rice[0][28] = 16'b10111_110111_11111;
        chicken_rice[0][29] = 16'b10111_110111_11111;
        chicken_rice[0][30] = 16'b10111_110111_11111;
        chicken_rice[0][31] = 16'b10111_110111_11111;
        chicken_rice[1][0] = 16'b10111_110111_11111;
        chicken_rice[1][1] = 16'b10111_110111_11111;
        chicken_rice[1][2] = 16'b10111_110111_11111;
        chicken_rice[1][3] = 16'b10111_110111_11111;
        chicken_rice[1][4] = 16'b10111_110111_11111;
        chicken_rice[1][5] = 16'b10111_110111_11111;
        chicken_rice[1][6] = 16'b10111_110111_11111;
        chicken_rice[1][7] = 16'b10111_110111_11111;
        chicken_rice[1][8] = 16'b10111_110111_11111;
        chicken_rice[1][9] = 16'b10111_110111_11111;
        chicken_rice[1][10] = 16'b10111_110111_11111;
        chicken_rice[1][11] = 16'b10111_110111_11111;
        chicken_rice[1][12] = 16'b10111_110111_11111;
        chicken_rice[1][13] = 16'b10111_110111_11111;
        chicken_rice[1][14] = 16'b10111_110111_11111;
        chicken_rice[1][15] = 16'b10111_110111_11111;
        chicken_rice[1][16] = 16'b10111_110111_11111;
        chicken_rice[1][17] = 16'b10111_110111_11111;
        chicken_rice[1][18] = 16'b10111_110111_11111;
        chicken_rice[1][19] = 16'b10111_110111_11111;
        chicken_rice[1][20] = 16'b10111_110111_11111;
        chicken_rice[1][21] = 16'b10111_110111_11111;
        chicken_rice[1][22] = 16'b10111_110111_11111;
        chicken_rice[1][23] = 16'b10111_110111_11111;
        chicken_rice[1][24] = 16'b10111_110111_11111;
        chicken_rice[1][25] = 16'b10111_110111_11111;
        chicken_rice[1][26] = 16'b10111_110111_11111;
        chicken_rice[1][27] = 16'b10111_110111_11111;
        chicken_rice[1][28] = 16'b10111_110111_11111;
        chicken_rice[1][29] = 16'b10111_110111_11111;
        chicken_rice[1][30] = 16'b10111_110111_11111;
        chicken_rice[1][31] = 16'b10111_110111_11111;
        chicken_rice[2][0] = 16'b10111_110111_11111;
        chicken_rice[2][1] = 16'b10111_110111_11111;
        chicken_rice[2][2] = 16'b10111_110111_11111;
        chicken_rice[2][3] = 16'b10111_110111_11111;
        chicken_rice[2][4] = 16'b10111_110111_11111;
        chicken_rice[2][5] = 16'b10111_110111_11111;
        chicken_rice[2][6] = 16'b10111_110111_11111;
        chicken_rice[2][7] = 16'b10111_110111_11111;
        chicken_rice[2][8] = 16'b10111_110111_11111;
        chicken_rice[2][9] = 16'b10111_110111_11111;
        chicken_rice[2][10] = 16'b10111_110111_11111;
        chicken_rice[2][11] = 16'b10111_110111_11111;
        chicken_rice[2][12] = 16'b10111_110111_11111;
        chicken_rice[2][13] = 16'b10111_110111_11111;
        chicken_rice[2][14] = 16'b10111_110111_11111;
        chicken_rice[2][15] = 16'b10111_110111_11111;
        chicken_rice[2][16] = 16'b10111_110111_11111;
        chicken_rice[2][17] = 16'b10111_110111_11111;
        chicken_rice[2][18] = 16'b10111_110111_11111;
        chicken_rice[2][19] = 16'b10111_110111_11111;
        chicken_rice[2][20] = 16'b10111_110111_11111;
        chicken_rice[2][21] = 16'b10111_110111_11111;
        chicken_rice[2][22] = 16'b10111_110111_11111;
        chicken_rice[2][23] = 16'b10111_110111_11111;
        chicken_rice[2][24] = 16'b10111_110111_11111;
        chicken_rice[2][25] = 16'b10111_110111_11111;
        chicken_rice[2][26] = 16'b10111_110111_11111;
        chicken_rice[2][27] = 16'b10111_110111_11111;
        chicken_rice[2][28] = 16'b10111_110111_11111;
        chicken_rice[2][29] = 16'b10111_110111_11111;
        chicken_rice[2][30] = 16'b10111_110111_11111;
        chicken_rice[2][31] = 16'b10111_110111_11111;
        chicken_rice[3][0] = 16'b10111_110111_11111;
        chicken_rice[3][1] = 16'b10111_110111_11111;
        chicken_rice[3][2] = 16'b10111_110111_11111;
        chicken_rice[3][3] = 16'b10111_110111_11111;
        chicken_rice[3][4] = 16'b10111_110111_11111;
        chicken_rice[3][5] = 16'b10111_110111_11111;
        chicken_rice[3][6] = 16'b10111_110111_11111;
        chicken_rice[3][7] = 16'b10111_110111_11111;
        chicken_rice[3][8] = 16'b10111_110111_11111;
        chicken_rice[3][9] = 16'b10111_110111_11111;
        chicken_rice[3][10] = 16'b10111_110111_11111;
        chicken_rice[3][11] = 16'b10111_110111_11111;
        chicken_rice[3][12] = 16'b10111_110111_11111;
        chicken_rice[3][13] = 16'b10111_110111_11111;
        chicken_rice[3][14] = 16'b10111_110111_11111;
        chicken_rice[3][15] = 16'b10111_110111_11111;
        chicken_rice[3][16] = 16'b10111_110111_11111;
        chicken_rice[3][17] = 16'b10111_110111_11111;
        chicken_rice[3][18] = 16'b10111_110111_11111;
        chicken_rice[3][19] = 16'b10111_110111_11111;
        chicken_rice[3][20] = 16'b10111_110111_11111;
        chicken_rice[3][21] = 16'b10111_110111_11111;
        chicken_rice[3][22] = 16'b10111_110111_11111;
        chicken_rice[3][23] = 16'b10111_110111_11111;
        chicken_rice[3][24] = 16'b10111_110111_11111;
        chicken_rice[3][25] = 16'b10111_110111_11111;
        chicken_rice[3][26] = 16'b10111_110111_11111;
        chicken_rice[3][27] = 16'b10111_110111_11111;
        chicken_rice[3][28] = 16'b10111_110111_11111;
        chicken_rice[3][29] = 16'b10111_110111_11111;
        chicken_rice[3][30] = 16'b10111_110111_11111;
        chicken_rice[3][31] = 16'b10111_110111_11111;
        chicken_rice[4][0] = 16'b10111_110111_11111;
        chicken_rice[4][1] = 16'b10111_110111_11111;
        chicken_rice[4][2] = 16'b10111_110111_11111;
        chicken_rice[4][3] = 16'b10111_110111_11111;
        chicken_rice[4][4] = 16'b10111_110111_11111;
        chicken_rice[4][5] = 16'b10111_110111_11111;
        chicken_rice[4][6] = 16'b10111_110111_11111;
        chicken_rice[4][7] = 16'b10111_110111_11111;
        chicken_rice[4][8] = 16'b10111_110111_11111;
        chicken_rice[4][9] = 16'b10111_110111_11111;
        chicken_rice[4][10] = 16'b10111_110111_11111;
        chicken_rice[4][11] = 16'b10111_110111_11111;
        chicken_rice[4][12] = 16'b10111_110111_11111;
        chicken_rice[4][13] = 16'b10111_110111_11111;
        chicken_rice[4][14] = 16'b10111_110111_11111;
        chicken_rice[4][15] = 16'b10111_110111_11111;
        chicken_rice[4][16] = 16'b10111_110111_11111;
        chicken_rice[4][17] = 16'b10111_110111_11111;
        chicken_rice[4][18] = 16'b10111_110111_11111;
        chicken_rice[4][19] = 16'b10111_110111_11111;
        chicken_rice[4][20] = 16'b10111_110111_11111;
        chicken_rice[4][21] = 16'b10111_110111_11111;
        chicken_rice[4][22] = 16'b10111_110111_11111;
        chicken_rice[4][23] = 16'b10111_110111_11111;
        chicken_rice[4][24] = 16'b10111_110111_11111;
        chicken_rice[4][25] = 16'b10111_110111_11111;
        chicken_rice[4][26] = 16'b10111_110111_11111;
        chicken_rice[4][27] = 16'b10111_110111_11111;
        chicken_rice[4][28] = 16'b10111_110111_11111;
        chicken_rice[4][29] = 16'b10111_110111_11111;
        chicken_rice[4][30] = 16'b10111_110111_11111;
        chicken_rice[4][31] = 16'b10111_110111_11111;
        chicken_rice[5][0] = 16'b10111_110111_11111;
        chicken_rice[5][1] = 16'b10111_110111_11111;
        chicken_rice[5][2] = 16'b10111_110111_11111;
        chicken_rice[5][3] = 16'b10111_110111_11111;
        chicken_rice[5][4] = 16'b10111_110111_11111;
        chicken_rice[5][5] = 16'b10111_110111_11111;
        chicken_rice[5][6] = 16'b10111_110111_11111;
        chicken_rice[5][7] = 16'b10111_110111_11111;
        chicken_rice[5][8] = 16'b10111_110111_11111;
        chicken_rice[5][9] = 16'b10111_110111_11111;
        chicken_rice[5][10] = 16'b10111_110111_11111;
        chicken_rice[5][11] = 16'b10111_110111_11111;
        chicken_rice[5][12] = 16'b11001_101001_01100;
        chicken_rice[5][13] = 16'b11010_101001_01100;
        chicken_rice[5][14] = 16'b11010_101010_01101;
        chicken_rice[5][15] = 16'b11010_101100_01110;
        chicken_rice[5][16] = 16'b11010_101011_01110;
        chicken_rice[5][17] = 16'b11100_110000_10000;
        chicken_rice[5][18] = 16'b11010_101100_01110;
        chicken_rice[5][19] = 16'b10111_110111_11111;
        chicken_rice[5][20] = 16'b10111_110111_11111;
        chicken_rice[5][21] = 16'b10111_110111_11111;
        chicken_rice[5][22] = 16'b10111_110111_11111;
        chicken_rice[5][23] = 16'b10111_110111_11111;
        chicken_rice[5][24] = 16'b10111_110111_11111;
        chicken_rice[5][25] = 16'b10111_110111_11111;
        chicken_rice[5][26] = 16'b10111_110111_11111;
        chicken_rice[5][27] = 16'b10111_110111_11111;
        chicken_rice[5][28] = 16'b10111_110111_11111;
        chicken_rice[5][29] = 16'b10111_110111_11111;
        chicken_rice[5][30] = 16'b10111_110111_11111;
        chicken_rice[5][31] = 16'b10111_110111_11111;
        chicken_rice[6][0] = 16'b10111_110111_11111;
        chicken_rice[6][1] = 16'b10111_110111_11111;
        chicken_rice[6][2] = 16'b10111_110111_11111;
        chicken_rice[6][3] = 16'b10111_110111_11111;
        chicken_rice[6][4] = 16'b10111_110111_11111;
        chicken_rice[6][5] = 16'b10111_110111_11111;
        chicken_rice[6][6] = 16'b10111_110111_11111;
        chicken_rice[6][7] = 16'b10111_110111_11111;
        chicken_rice[6][8] = 16'b10111_110111_11111;
        chicken_rice[6][9] = 16'b11001_101000_01100;
        chicken_rice[6][10] = 16'b11100_101111_10000;
        chicken_rice[6][11] = 16'b11011_101111_01111;
        chicken_rice[6][12] = 16'b11011_101101_01111;
        chicken_rice[6][13] = 16'b11011_101110_01111;
        chicken_rice[6][14] = 16'b11100_101111_10000;
        chicken_rice[6][15] = 16'b11100_110000_10000;
        chicken_rice[6][16] = 16'b11100_101111_10000;
        chicken_rice[6][17] = 16'b11100_110001_10001;
        chicken_rice[6][18] = 16'b11100_110000_10000;
        chicken_rice[6][19] = 16'b11100_110001_10001;
        chicken_rice[6][20] = 16'b11100_110001_10001;
        chicken_rice[6][21] = 16'b11100_110000_10000;
        chicken_rice[6][22] = 16'b11010_101100_01110;
        chicken_rice[6][23] = 16'b10111_110111_11111;
        chicken_rice[6][24] = 16'b10111_110111_11111;
        chicken_rice[6][25] = 16'b10111_110111_11111;
        chicken_rice[6][26] = 16'b10111_110111_11111;
        chicken_rice[6][27] = 16'b10111_110111_11111;
        chicken_rice[6][28] = 16'b10111_110111_11111;
        chicken_rice[6][29] = 16'b10111_110111_11111;
        chicken_rice[6][30] = 16'b10111_110111_11111;
        chicken_rice[6][31] = 16'b10111_110111_11111;
        chicken_rice[7][0] = 16'b10111_110111_11111;
        chicken_rice[7][1] = 16'b10111_110111_11111;
        chicken_rice[7][2] = 16'b10111_110111_11111;
        chicken_rice[7][3] = 16'b10111_110111_11111;
        chicken_rice[7][4] = 16'b10111_110111_11111;
        chicken_rice[7][5] = 16'b10111_110111_11111;
        chicken_rice[7][6] = 16'b10111_110111_11111;
        chicken_rice[7][7] = 16'b11001_101000_01100;
        chicken_rice[7][8] = 16'b11100_101111_01111;
        chicken_rice[7][9] = 16'b11011_101110_01111;
        chicken_rice[7][10] = 16'b11011_101101_01111;
        chicken_rice[7][11] = 16'b11011_101110_01111;
        chicken_rice[7][12] = 16'b11010_101011_01110;
        chicken_rice[7][13] = 16'b11010_101101_01111;
        chicken_rice[7][14] = 16'b11011_101110_01111;
        chicken_rice[7][15] = 16'b11011_101110_01111;
        chicken_rice[7][16] = 16'b11011_101110_01111;
        chicken_rice[7][17] = 16'b11011_101111_10000;
        chicken_rice[7][18] = 16'b11100_110000_10000;
        chicken_rice[7][19] = 16'b11100_110000_10000;
        chicken_rice[7][20] = 16'b11100_110000_10000;
        chicken_rice[7][21] = 16'b11100_110000_10001;
        chicken_rice[7][22] = 16'b11100_110000_10000;
        chicken_rice[7][23] = 16'b11100_110001_10001;
        chicken_rice[7][24] = 16'b10111_110111_11111;
        chicken_rice[7][25] = 16'b10111_110111_11111;
        chicken_rice[7][26] = 16'b10111_110111_11111;
        chicken_rice[7][27] = 16'b10111_110111_11111;
        chicken_rice[7][28] = 16'b10111_110111_11111;
        chicken_rice[7][29] = 16'b10111_110111_11111;
        chicken_rice[7][30] = 16'b10111_110111_11111;
        chicken_rice[7][31] = 16'b10111_110111_11111;
        chicken_rice[8][0] = 16'b10111_110111_11111;
        chicken_rice[8][1] = 16'b10111_110111_11111;
        chicken_rice[8][2] = 16'b10111_110111_11111;
        chicken_rice[8][3] = 16'b10111_110111_11111;
        chicken_rice[8][4] = 16'b10111_110111_11111;
        chicken_rice[8][5] = 16'b10111_110111_11111;
        chicken_rice[8][6] = 16'b11001_101000_01100;
        chicken_rice[8][7] = 16'b11011_101111_10000;
        chicken_rice[8][8] = 16'b11011_101101_01110;
        chicken_rice[8][9] = 16'b10110_011111_00111;
        chicken_rice[8][10] = 16'b10110_011110_00110;
        chicken_rice[8][11] = 16'b11000_100011_01000;
        chicken_rice[8][12] = 16'b11000_100001_00110;
        chicken_rice[8][13] = 16'b11000_100001_00111;
        chicken_rice[8][14] = 16'b11000_100010_00111;
        chicken_rice[8][15] = 16'b10110_011101_00101;
        chicken_rice[8][16] = 16'b11000_100100_01001;
        chicken_rice[8][17] = 16'b11001_100111_01011;
        chicken_rice[8][18] = 16'b11000_100110_01011;
        chicken_rice[8][19] = 16'b11001_101001_01100;
        chicken_rice[8][20] = 16'b11010_101010_01101;
        chicken_rice[8][21] = 16'b11010_101011_01101;
        chicken_rice[8][22] = 16'b11011_101111_10000;
        chicken_rice[8][23] = 16'b11100_110001_10000;
        chicken_rice[8][24] = 16'b11100_110001_10001;
        chicken_rice[8][25] = 16'b11010_101010_01101;
        chicken_rice[8][26] = 16'b10111_110111_11111;
        chicken_rice[8][27] = 16'b10111_110111_11111;
        chicken_rice[8][28] = 16'b10111_110111_11111;
        chicken_rice[8][29] = 16'b10111_110111_11111;
        chicken_rice[8][30] = 16'b10111_110111_11111;
        chicken_rice[8][31] = 16'b10111_110111_11111;
        chicken_rice[9][0] = 16'b10111_110111_11111;
        chicken_rice[9][1] = 16'b10111_110111_11111;
        chicken_rice[9][2] = 16'b10111_110111_11111;
        chicken_rice[9][3] = 16'b10111_110111_11111;
        chicken_rice[9][4] = 16'b11001_101010_01110;
        chicken_rice[9][5] = 16'b11100_110000_10000;
        chicken_rice[9][6] = 16'b11100_110000_10000;
        chicken_rice[9][7] = 16'b11001_101000_01100;
        chicken_rice[9][8] = 16'b10111_011110_00101;
        chicken_rice[9][9] = 16'b10111_011010_00011;
        chicken_rice[9][10] = 16'b11001_011110_00011;
        chicken_rice[9][11] = 16'b11011_100110_00111;
        chicken_rice[9][12] = 16'b11100_101100_01101;
        chicken_rice[9][13] = 16'b11101_110000_10000;
        chicken_rice[9][14] = 16'b11011_101000_01010;
        chicken_rice[9][15] = 16'b11000_100000_00101;
        chicken_rice[9][16] = 16'b10110_011011_00100;
        chicken_rice[9][17] = 16'b10111_100001_00111;
        chicken_rice[9][18] = 16'b11000_100011_01000;
        chicken_rice[9][19] = 16'b11001_101001_01100;
        chicken_rice[9][20] = 16'b11000_100110_01011;
        chicken_rice[9][21] = 16'b11000_100110_01010;
        chicken_rice[9][22] = 16'b11000_100011_01001;
        chicken_rice[9][23] = 16'b11000_100011_01001;
        chicken_rice[9][24] = 16'b11100_101111_10000;
        chicken_rice[9][25] = 16'b11011_101111_10000;
        chicken_rice[9][26] = 16'b11100_101111_10000;
        chicken_rice[9][27] = 16'b11001_101010_01101;
        chicken_rice[9][28] = 16'b10111_110111_11111;
        chicken_rice[9][29] = 16'b10111_110111_11111;
        chicken_rice[9][30] = 16'b10111_110111_11111;
        chicken_rice[9][31] = 16'b10111_110111_11111;
        chicken_rice[10][0] = 16'b10111_110111_11111;
        chicken_rice[10][1] = 16'b10111_110111_11111;
        chicken_rice[10][2] = 16'b10111_110111_11111;
        chicken_rice[10][3] = 16'b11011_101111_10000;
        chicken_rice[10][4] = 16'b11100_110000_10001;
        chicken_rice[10][5] = 16'b11100_110000_10000;
        chicken_rice[10][6] = 16'b11010_101010_01101;
        chicken_rice[10][7] = 16'b11000_100001_00111;
        chicken_rice[10][8] = 16'b10111_011011_00010;
        chicken_rice[10][9] = 16'b11011_100000_00010;
        chicken_rice[10][10] = 16'b11011_100000_00010;
        chicken_rice[10][11] = 16'b11010_100010_00100;
        chicken_rice[10][12] = 16'b11010_100001_00100;
        chicken_rice[10][13] = 16'b11011_100111_01001;
        chicken_rice[10][14] = 16'b11100_101010_01011;
        chicken_rice[10][15] = 16'b11011_101000_01010;
        chicken_rice[10][16] = 16'b11001_011111_00100;
        chicken_rice[10][17] = 16'b11001_100101_01001;
        chicken_rice[10][18] = 16'b11010_101000_01011;
        chicken_rice[10][19] = 16'b11100_110001_10001;
        chicken_rice[10][20] = 16'b11010_101011_01101;
        chicken_rice[10][21] = 16'b11010_101010_01101;
        chicken_rice[10][22] = 16'b11011_101101_01110;
        chicken_rice[10][23] = 16'b11011_101100_01110;
        chicken_rice[10][24] = 16'b11000_100100_01001;
        chicken_rice[10][25] = 16'b11010_101011_01101;
        chicken_rice[10][26] = 16'b11100_101111_10000;
        chicken_rice[10][27] = 16'b11100_110000_10000;
        chicken_rice[10][28] = 16'b11010_101100_01110;
        chicken_rice[10][29] = 16'b10111_110111_11111;
        chicken_rice[10][30] = 16'b10111_110111_11111;
        chicken_rice[10][31] = 16'b10111_110111_11111;
        chicken_rice[11][0] = 16'b10111_110111_11111;
        chicken_rice[11][1] = 16'b10111_110111_11111;
        chicken_rice[11][2] = 16'b10111_110111_11111;
        chicken_rice[11][3] = 16'b11100_110001_10001;
        chicken_rice[11][4] = 16'b11100_110001_10001;
        chicken_rice[11][5] = 16'b11100_110000_10000;
        chicken_rice[11][6] = 16'b11000_100011_01001;
        chicken_rice[11][7] = 16'b10111_011010_00010;
        chicken_rice[11][8] = 16'b11000_011011_00001;
        chicken_rice[11][9] = 16'b11100_100101_00100;
        chicken_rice[11][10] = 16'b11100_100101_00100;
        chicken_rice[11][11] = 16'b11100_100110_00101;
        chicken_rice[11][12] = 16'b11101_100111_00110;
        chicken_rice[11][13] = 16'b11100_101001_01000;
        chicken_rice[11][14] = 16'b11001_100011_00111;
        chicken_rice[11][15] = 16'b11011_101001_01011;
        chicken_rice[11][16] = 16'b11010_100110_01001;
        chicken_rice[11][17] = 16'b11000_100010_01000;
        chicken_rice[11][18] = 16'b11011_101110_01111;
        chicken_rice[11][19] = 16'b11100_110001_10001;
        chicken_rice[11][20] = 16'b11100_110000_10000;
        chicken_rice[11][21] = 16'b11011_101111_01111;
        chicken_rice[11][22] = 16'b11100_110001_10001;
        chicken_rice[11][23] = 16'b11100_110010_10001;
        chicken_rice[11][24] = 16'b11011_101101_01110;
        chicken_rice[11][25] = 16'b10111_100010_01001;
        chicken_rice[11][26] = 16'b11010_101011_01110;
        chicken_rice[11][27] = 16'b11011_101111_10000;
        chicken_rice[11][28] = 16'b11100_110000_10001;
        chicken_rice[11][29] = 16'b10111_110111_11111;
        chicken_rice[11][30] = 16'b10111_110111_11111;
        chicken_rice[11][31] = 16'b10111_110111_11111;
        chicken_rice[12][0] = 16'b10111_110111_11111;
        chicken_rice[12][1] = 16'b10111_110111_11111;
        chicken_rice[12][2] = 16'b11011_101111_10000;
        chicken_rice[12][3] = 16'b11100_110000_10001;
        chicken_rice[12][4] = 16'b11100_110000_10000;
        chicken_rice[12][5] = 16'b11010_101001_01100;
        chicken_rice[12][6] = 16'b11000_011101_00100;
        chicken_rice[12][7] = 16'b11010_011101_00001;
        chicken_rice[12][8] = 16'b11001_011100_00000;
        chicken_rice[12][9] = 16'b11000_011000_00000;
        chicken_rice[12][10] = 16'b11100_100110_00101;
        chicken_rice[12][11] = 16'b11100_101001_01000;
        chicken_rice[12][12] = 16'b11101_101101_01011;
        chicken_rice[12][13] = 16'b11100_101010_01001;
        chicken_rice[12][14] = 16'b11011_100110_00111;
        chicken_rice[12][15] = 16'b11010_100100_00110;
        chicken_rice[12][16] = 16'b11010_100001_00100;
        chicken_rice[12][17] = 16'b10111_011111_00111;
        chicken_rice[12][18] = 16'b11010_101100_01101;
        chicken_rice[12][19] = 16'b11100_110000_10000;
        chicken_rice[12][20] = 16'b11101_110011_10010;
        chicken_rice[12][21] = 16'b11011_101111_10000;
        chicken_rice[12][22] = 16'b11011_101111_10000;
        chicken_rice[12][23] = 16'b11101_110011_10010;
        chicken_rice[12][24] = 16'b11100_110010_10001;
        chicken_rice[12][25] = 16'b11010_101010_01101;
        chicken_rice[12][26] = 16'b11000_100011_01001;
        chicken_rice[12][27] = 16'b11011_101110_01111;
        chicken_rice[12][28] = 16'b11100_110001_10001;
        chicken_rice[12][29] = 16'b11100_110001_10001;
        chicken_rice[12][30] = 16'b10111_110111_11111;
        chicken_rice[12][31] = 16'b10111_110111_11111;
        chicken_rice[13][0] = 16'b10111_110111_11111;
        chicken_rice[13][1] = 16'b10111_110111_11111;
        chicken_rice[13][2] = 16'b11100_110010_10010;
        chicken_rice[13][3] = 16'b11100_110001_10001;
        chicken_rice[13][4] = 16'b11100_110000_10000;
        chicken_rice[13][5] = 16'b11001_101000_01011;
        chicken_rice[13][6] = 16'b10111_011001_00001;
        chicken_rice[13][7] = 16'b11010_100001_00011;
        chicken_rice[13][8] = 16'b11011_100010_00011;
        chicken_rice[13][9] = 16'b10110_010110_00000;
        chicken_rice[13][10] = 16'b10111_011000_00000;
        chicken_rice[13][11] = 16'b11011_100010_00011;
        chicken_rice[13][12] = 16'b11011_100100_00100;
        chicken_rice[13][13] = 16'b11100_101011_01010;
        chicken_rice[13][14] = 16'b11011_100101_00101;
        chicken_rice[13][15] = 16'b11010_100010_00100;
        chicken_rice[13][16] = 16'b11010_011110_00010;
        chicken_rice[13][17] = 16'b11000_011011_00001;
        chicken_rice[13][18] = 16'b11100_101111_10000;
        chicken_rice[13][19] = 16'b11101_110011_10010;
        chicken_rice[13][20] = 16'b11100_110000_10000;
        chicken_rice[13][21] = 16'b11011_101111_10000;
        chicken_rice[13][22] = 16'b11101_110011_10010;
        chicken_rice[13][23] = 16'b11101_110100_10010;
        chicken_rice[13][24] = 16'b11100_110010_10001;
        chicken_rice[13][25] = 16'b11100_110000_10001;
        chicken_rice[13][26] = 16'b11001_100110_01010;
        chicken_rice[13][27] = 16'b11010_101100_01110;
        chicken_rice[13][28] = 16'b11100_110000_10000;
        chicken_rice[13][29] = 16'b11100_110010_10001;
        chicken_rice[13][30] = 16'b10111_110111_11111;
        chicken_rice[13][31] = 16'b10111_110111_11111;
        chicken_rice[14][0] = 16'b10111_110111_11111;
        chicken_rice[14][1] = 16'b10111_110111_11111;
        chicken_rice[14][2] = 16'b11100_110010_10010;
        chicken_rice[14][3] = 16'b11100_110001_10001;
        chicken_rice[14][4] = 16'b11011_101110_01111;
        chicken_rice[14][5] = 16'b10110_011001_00010;
        chicken_rice[14][6] = 16'b10101_010110_00001;
        chicken_rice[14][7] = 16'b10111_011001_00001;
        chicken_rice[14][8] = 16'b11011_100010_00011;
        chicken_rice[14][9] = 16'b11100_100110_00100;
        chicken_rice[14][10] = 16'b11100_100101_00100;
        chicken_rice[14][11] = 16'b11001_011101_00001;
        chicken_rice[14][12] = 16'b11001_011110_00001;
        chicken_rice[14][13] = 16'b11010_100010_00100;
        chicken_rice[14][14] = 16'b11100_101000_00111;
        chicken_rice[14][15] = 16'b11100_100110_00110;
        chicken_rice[14][16] = 16'b11100_100110_00110;
        chicken_rice[14][17] = 16'b11010_100010_00100;
        chicken_rice[14][18] = 16'b11010_101011_01110;
        chicken_rice[14][19] = 16'b11100_110001_10001;
        chicken_rice[14][20] = 16'b11100_110001_10001;
        chicken_rice[14][21] = 16'b11100_110001_10001;
        chicken_rice[14][22] = 16'b11101_110100_10011;
        chicken_rice[14][23] = 16'b11100_110010_10010;
        chicken_rice[14][24] = 16'b11101_110101_10011;
        chicken_rice[14][25] = 16'b11100_110010_10010;
        chicken_rice[14][26] = 16'b11011_101110_01111;
        chicken_rice[14][27] = 16'b11001_100111_01011;
        chicken_rice[14][28] = 16'b11100_110000_10000;
        chicken_rice[14][29] = 16'b11100_110001_10001;
        chicken_rice[14][30] = 16'b10111_110111_11111;
        chicken_rice[14][31] = 16'b10111_110111_11111;
        chicken_rice[15][0] = 16'b10111_110111_11111;
        chicken_rice[15][1] = 16'b10111_110111_11111;
        chicken_rice[15][2] = 16'b11100_110011_10010;
        chicken_rice[15][3] = 16'b11100_110010_10001;
        chicken_rice[15][4] = 16'b11010_101100_01110;
        chicken_rice[15][5] = 16'b10110_011000_00001;
        chicken_rice[15][6] = 16'b11010_011110_00001;
        chicken_rice[15][7] = 16'b10110_010110_00000;
        chicken_rice[15][8] = 16'b11001_011101_00010;
        chicken_rice[15][9] = 16'b11101_101010_00111;
        chicken_rice[15][10] = 16'b11101_101110_01011;
        chicken_rice[15][11] = 16'b11100_101001_01000;
        chicken_rice[15][12] = 16'b11100_100111_00111;
        chicken_rice[15][13] = 16'b11010_100010_00101;
        chicken_rice[15][14] = 16'b11010_100010_00101;
        chicken_rice[15][15] = 16'b11000_011100_00010;
        chicken_rice[15][16] = 16'b11000_011100_00010;
        chicken_rice[15][17] = 16'b11010_100010_00101;
        chicken_rice[15][18] = 16'b11011_101110_01111;
        chicken_rice[15][19] = 16'b11100_110010_10010;
        chicken_rice[15][20] = 16'b11101_110101_10100;
        chicken_rice[15][21] = 16'b11101_110011_10010;
        chicken_rice[15][22] = 16'b11101_110100_10011;
        chicken_rice[15][23] = 16'b11101_110110_10100;
        chicken_rice[15][24] = 16'b11100_110011_10010;
        chicken_rice[15][25] = 16'b11101_110100_10011;
        chicken_rice[15][26] = 16'b11100_110000_10000;
        chicken_rice[15][27] = 16'b11001_100111_01011;
        chicken_rice[15][28] = 16'b11100_110000_10000;
        chicken_rice[15][29] = 16'b11100_110010_10001;
        chicken_rice[15][30] = 16'b10111_110111_11111;
        chicken_rice[15][31] = 16'b10111_110111_11111;
        chicken_rice[16][0] = 16'b10111_110111_11111;
        chicken_rice[16][1] = 16'b10111_110111_11111;
        chicken_rice[16][2] = 16'b11100_110010_10010;
        chicken_rice[16][3] = 16'b11100_110001_10001;
        chicken_rice[16][4] = 16'b11010_101011_01101;
        chicken_rice[16][5] = 16'b10111_011001_00010;
        chicken_rice[16][6] = 16'b11010_100000_00010;
        chicken_rice[16][7] = 16'b11011_100100_00100;
        chicken_rice[16][8] = 16'b11010_011110_00001;
        chicken_rice[16][9] = 16'b11011_100000_00001;
        chicken_rice[16][10] = 16'b11101_101001_00111;
        chicken_rice[16][11] = 16'b11101_110000_01111;
        chicken_rice[16][12] = 16'b11101_110000_01111;
        chicken_rice[16][13] = 16'b11100_101010_01001;
        chicken_rice[16][14] = 16'b11011_100110_00111;
        chicken_rice[16][15] = 16'b11001_011110_00001;
        chicken_rice[16][16] = 16'b11001_011011_00000;
        chicken_rice[16][17] = 16'b11100_100111_00111;
        chicken_rice[16][18] = 16'b11100_110011_10010;
        chicken_rice[16][19] = 16'b11101_110100_10011;
        chicken_rice[16][20] = 16'b11101_110110_10100;
        chicken_rice[16][21] = 16'b11100_110011_10010;
        chicken_rice[16][22] = 16'b11100_110010_10010;
        chicken_rice[16][23] = 16'b11110_110110_10101;
        chicken_rice[16][24] = 16'b11101_110011_10011;
        chicken_rice[16][25] = 16'b11101_110011_10011;
        chicken_rice[16][26] = 16'b11100_110001_10001;
        chicken_rice[16][27] = 16'b11001_101000_01011;
        chicken_rice[16][28] = 16'b11100_110000_10000;
        chicken_rice[16][29] = 16'b11100_110001_10001;
        chicken_rice[16][30] = 16'b10111_110111_11111;
        chicken_rice[16][31] = 16'b10111_110111_11111;
        chicken_rice[17][0] = 16'b10111_110111_11111;
        chicken_rice[17][1] = 16'b10111_110111_11111;
        chicken_rice[17][2] = 16'b11100_110010_10010;
        chicken_rice[17][3] = 16'b11100_110001_10001;
        chicken_rice[17][4] = 16'b11011_101110_01111;
        chicken_rice[17][5] = 16'b10111_011010_00001;
        chicken_rice[17][6] = 16'b11011_100001_00011;
        chicken_rice[17][7] = 16'b11100_100111_00111;
        chicken_rice[17][8] = 16'b11100_100111_00110;
        chicken_rice[17][9] = 16'b11011_100000_00001;
        chicken_rice[17][10] = 16'b11010_011101_00000;
        chicken_rice[17][11] = 16'b11010_100000_00011;
        chicken_rice[17][12] = 16'b11011_100011_00101;
        chicken_rice[17][13] = 16'b11011_100101_00110;
        chicken_rice[17][14] = 16'b11011_100110_00111;
        chicken_rice[17][15] = 16'b11001_011100_00001;
        chicken_rice[17][16] = 16'b10111_010111_00000;
        chicken_rice[17][17] = 16'b11100_101000_00111;
        chicken_rice[17][18] = 16'b11101_110100_10011;
        chicken_rice[17][19] = 16'b11110_110110_10101;
        chicken_rice[17][20] = 16'b11101_110100_10011;
        chicken_rice[17][21] = 16'b11110_110110_10101;
        chicken_rice[17][22] = 16'b11101_110011_10011;
        chicken_rice[17][23] = 16'b11100_110011_10010;
        chicken_rice[17][24] = 16'b11101_110110_10100;
        chicken_rice[17][25] = 16'b11101_110011_10010;
        chicken_rice[17][26] = 16'b11011_101111_10000;
        chicken_rice[17][27] = 16'b11001_101001_01100;
        chicken_rice[17][28] = 16'b11011_110000_10000;
        chicken_rice[17][29] = 16'b11100_110001_10001;
        chicken_rice[17][30] = 16'b10111_110111_11111;
        chicken_rice[17][31] = 16'b10111_110111_11111;
        chicken_rice[18][0] = 16'b10111_110111_11111;
        chicken_rice[18][1] = 16'b10111_110111_11111;
        chicken_rice[18][2] = 16'b11100_110010_10010;
        chicken_rice[18][3] = 16'b11100_110010_10001;
        chicken_rice[18][4] = 16'b11100_110000_10000;
        chicken_rice[18][5] = 16'b11010_101001_01011;
        chicken_rice[18][6] = 16'b11000_011001_00000;
        chicken_rice[18][7] = 16'b11001_011111_00010;
        chicken_rice[18][8] = 16'b11100_101000_00111;
        chicken_rice[18][9] = 16'b11101_101011_01010;
        chicken_rice[18][10] = 16'b11100_101011_01001;
        chicken_rice[18][11] = 16'b11011_100011_00101;
        chicken_rice[18][12] = 16'b11001_011110_00011;
        chicken_rice[18][13] = 16'b11010_100000_00011;
        chicken_rice[18][14] = 16'b10111_011001_00000;
        chicken_rice[18][15] = 16'b10111_011001_00000;
        chicken_rice[18][16] = 16'b11000_011010_00000;
        chicken_rice[18][17] = 16'b11100_110010_10010;
        chicken_rice[18][18] = 16'b11101_110110_10100;
        chicken_rice[18][19] = 16'b11101_110100_10011;
        chicken_rice[18][20] = 16'b11101_110100_10011;
        chicken_rice[18][21] = 16'b11101_110110_10101;
        chicken_rice[18][22] = 16'b11101_110111_10101;
        chicken_rice[18][23] = 16'b11101_110100_10011;
        chicken_rice[18][24] = 16'b11101_110100_10011;
        chicken_rice[18][25] = 16'b11101_110011_10011;
        chicken_rice[18][26] = 16'b11010_101011_01101;
        chicken_rice[18][27] = 16'b11011_101110_01111;
        chicken_rice[18][28] = 16'b11100_110000_10000;
        chicken_rice[18][29] = 16'b11100_110000_10000;
        chicken_rice[18][30] = 16'b10111_110111_11111;
        chicken_rice[18][31] = 16'b10111_110111_11111;
        chicken_rice[19][0] = 16'b10111_110111_11111;
        chicken_rice[19][1] = 16'b10111_110111_11111;
        chicken_rice[19][2] = 16'b10111_110111_11111;
        chicken_rice[19][3] = 16'b11100_110010_10010;
        chicken_rice[19][4] = 16'b11100_110000_10000;
        chicken_rice[19][5] = 16'b11100_110000_10000;
        chicken_rice[19][6] = 16'b11011_100010_00100;
        chicken_rice[19][7] = 16'b11001_011110_00010;
        chicken_rice[19][8] = 16'b11001_100000_00011;
        chicken_rice[19][9] = 16'b11100_101000_01000;
        chicken_rice[19][10] = 16'b11100_101011_01010;
        chicken_rice[19][11] = 16'b11100_101010_01001;
        chicken_rice[19][12] = 16'b11100_101010_01001;
        chicken_rice[19][13] = 16'b11010_100010_00100;
        chicken_rice[19][14] = 16'b11010_100010_00100;
        chicken_rice[19][15] = 16'b11001_011110_00010;
        chicken_rice[19][16] = 16'b11011_100100_00101;
        chicken_rice[19][17] = 16'b11101_110100_10100;
        chicken_rice[19][18] = 16'b11101_110100_10011;
        chicken_rice[19][19] = 16'b11101_110110_10101;
        chicken_rice[19][20] = 16'b11101_110100_10011;
        chicken_rice[19][21] = 16'b11101_110100_10011;
        chicken_rice[19][22] = 16'b11101_110110_10101;
        chicken_rice[19][23] = 16'b11101_110110_10100;
        chicken_rice[19][24] = 16'b11101_110101_10100;
        chicken_rice[19][25] = 16'b11100_110001_10001;
        chicken_rice[19][26] = 16'b11011_101110_01111;
        chicken_rice[19][27] = 16'b11011_101110_01111;
        chicken_rice[19][28] = 16'b11100_110000_10000;
        chicken_rice[19][29] = 16'b10111_110111_11111;
        chicken_rice[19][30] = 16'b10111_110111_11111;
        chicken_rice[19][31] = 16'b10111_110111_11111;
        chicken_rice[20][0] = 16'b10111_110111_11111;
        chicken_rice[20][1] = 16'b10111_110111_11111;
        chicken_rice[20][2] = 16'b10111_110111_11111;
        chicken_rice[20][3] = 16'b11100_110001_10001;
        chicken_rice[20][4] = 16'b11100_110001_10001;
        chicken_rice[20][5] = 16'b11100_110000_10001;
        chicken_rice[20][6] = 16'b11100_101111_01111;
        chicken_rice[20][7] = 16'b11011_100001_00011;
        chicken_rice[20][8] = 16'b11011_100010_00011;
        chicken_rice[20][9] = 16'b11010_100001_00011;
        chicken_rice[20][10] = 16'b11011_100001_00011;
        chicken_rice[20][11] = 16'b11011_100101_00101;
        chicken_rice[20][12] = 16'b11011_100100_00101;
        chicken_rice[20][13] = 16'b11010_100010_00100;
        chicken_rice[20][14] = 16'b11000_011100_00001;
        chicken_rice[20][15] = 16'b11001_011100_00001;
        chicken_rice[20][16] = 16'b11100_110010_10010;
        chicken_rice[20][17] = 16'b11110_110110_10101;
        chicken_rice[20][18] = 16'b11101_110100_10011;
        chicken_rice[20][19] = 16'b11110_110111_10101;
        chicken_rice[20][20] = 16'b11110_110111_10101;
        chicken_rice[20][21] = 16'b11101_110100_10011;
        chicken_rice[20][22] = 16'b11101_110101_10100;
        chicken_rice[20][23] = 16'b11101_110100_10011;
        chicken_rice[20][24] = 16'b11100_110011_10010;
        chicken_rice[20][25] = 16'b10010_100100_01010;
        chicken_rice[20][26] = 16'b11010_101101_01111;
        chicken_rice[20][27] = 16'b11011_101110_01111;
        chicken_rice[20][28] = 16'b11011_110000_10000;
        chicken_rice[20][29] = 16'b10111_110111_11111;
        chicken_rice[20][30] = 16'b10111_110111_11111;
        chicken_rice[20][31] = 16'b10111_110111_11111;
        chicken_rice[21][0] = 16'b10111_110111_11111;
        chicken_rice[21][1] = 16'b10111_110111_11111;
        chicken_rice[21][2] = 16'b10111_110111_11111;
        chicken_rice[21][3] = 16'b10111_110111_11111;
        chicken_rice[21][4] = 16'b11011_101111_10000;
        chicken_rice[21][5] = 16'b11100_110001_10001;
        chicken_rice[21][6] = 16'b11100_110001_10001;
        chicken_rice[21][7] = 16'b11010_100111_01010;
        chicken_rice[21][8] = 16'b11011_100011_00100;
        chicken_rice[21][9] = 16'b11100_101010_01001;
        chicken_rice[21][10] = 16'b11100_100100_00100;
        chicken_rice[21][11] = 16'b11010_100000_00011;
        chicken_rice[21][12] = 16'b11000_011100_00010;
        chicken_rice[21][13] = 16'b10111_011010_00001;
        chicken_rice[21][14] = 16'b11000_011011_00001;
        chicken_rice[21][15] = 16'b11010_101001_01100;
        chicken_rice[21][16] = 16'b11110_110110_10101;
        chicken_rice[21][17] = 16'b11110_111000_10110;
        chicken_rice[21][18] = 16'b11110_111000_10110;
        chicken_rice[21][19] = 16'b11110_110111_10101;
        chicken_rice[21][20] = 16'b11101_110110_10100;
        chicken_rice[21][21] = 16'b11110_110111_10101;
        chicken_rice[21][22] = 16'b11110_110110_10101;
        chicken_rice[21][23] = 16'b11101_110110_10100;
        chicken_rice[21][24] = 16'b10010_100100_01010;
        chicken_rice[21][25] = 16'b01101_011011_00101;
        chicken_rice[21][26] = 16'b11010_101100_01110;
        chicken_rice[21][27] = 16'b11011_101110_01111;
        chicken_rice[21][28] = 16'b10111_110111_11111;
        chicken_rice[21][29] = 16'b10111_110111_11111;
        chicken_rice[21][30] = 16'b10111_110111_11111;
        chicken_rice[21][31] = 16'b10111_110111_11111;
        chicken_rice[22][0] = 16'b10111_110111_11111;
        chicken_rice[22][1] = 16'b10111_110111_11111;
        chicken_rice[22][2] = 16'b10111_110111_11111;
        chicken_rice[22][3] = 16'b10111_110111_11111;
        chicken_rice[22][4] = 16'b10111_110111_11111;
        chicken_rice[22][5] = 16'b11011_101110_01111;
        chicken_rice[22][6] = 16'b11011_101110_01111;
        chicken_rice[22][7] = 16'b11011_101101_01110;
        chicken_rice[22][8] = 16'b11010_100110_01000;
        chicken_rice[22][9] = 16'b11100_100111_00110;
        chicken_rice[22][10] = 16'b11101_101110_01100;
        chicken_rice[22][11] = 16'b11101_101101_01011;
        chicken_rice[22][12] = 16'b11010_100101_01000;
        chicken_rice[22][13] = 16'b11010_100110_01001;
        chicken_rice[22][14] = 16'b11000_011101_00001;
        chicken_rice[22][15] = 16'b11000_100011_01000;
        chicken_rice[22][16] = 16'b11110_111000_10110;
        chicken_rice[22][17] = 16'b11110_111000_10110;
        chicken_rice[22][18] = 16'b11110_110111_10101;
        chicken_rice[22][19] = 16'b11110_110111_10101;
        chicken_rice[22][20] = 16'b11101_110101_10100;
        chicken_rice[22][21] = 16'b11101_110111_10101;
        chicken_rice[22][22] = 16'b11110_111000_10110;
        chicken_rice[22][23] = 16'b11101_110110_10100;
        chicken_rice[22][24] = 16'b01110_011110_00111;
        chicken_rice[22][25] = 16'b01100_011010_00101;
        chicken_rice[22][26] = 16'b11001_101011_01110;
        chicken_rice[22][27] = 16'b10111_110111_11111;
        chicken_rice[22][28] = 16'b10111_110111_11111;
        chicken_rice[22][29] = 16'b10111_110111_11111;
        chicken_rice[22][30] = 16'b10111_110111_11111;
        chicken_rice[22][31] = 16'b10111_110111_11111;
        chicken_rice[23][0] = 16'b10111_110111_11111;
        chicken_rice[23][1] = 16'b10111_110111_11111;
        chicken_rice[23][2] = 16'b10111_110111_11111;
        chicken_rice[23][3] = 16'b10111_110111_11111;
        chicken_rice[23][4] = 16'b10111_110111_11111;
        chicken_rice[23][5] = 16'b10111_110111_11111;
        chicken_rice[23][6] = 16'b10111_110111_11111;
        chicken_rice[23][7] = 16'b10111_110111_11111;
        chicken_rice[23][8] = 16'b11100_110000_10000;
        chicken_rice[23][9] = 16'b11100_110001_10001;
        chicken_rice[23][10] = 16'b11100_110001_10001;
        chicken_rice[23][11] = 16'b11100_110000_10000;
        chicken_rice[23][12] = 16'b11100_110000_10000;
        chicken_rice[23][13] = 16'b11100_110000_10000;
        chicken_rice[23][14] = 16'b11011_101101_01110;
        chicken_rice[23][15] = 16'b11011_101101_01110;
        chicken_rice[23][16] = 16'b10001_100010_01001;
        chicken_rice[23][17] = 16'b10010_100100_01010;
        chicken_rice[23][18] = 16'b10010_100100_01010;
        chicken_rice[23][19] = 16'b10001_100010_01001;
        chicken_rice[23][20] = 16'b01111_011111_01000;
        chicken_rice[23][21] = 16'b10100_100111_01011;
        chicken_rice[23][22] = 16'b10001_100011_01001;
        chicken_rice[23][23] = 16'b10100_100111_01011;
        chicken_rice[23][24] = 16'b01101_011100_00110;
        chicken_rice[23][25] = 16'b01101_011011_00101;
        chicken_rice[23][26] = 16'b10111_110111_11111;
        chicken_rice[23][27] = 16'b10111_110111_11111;
        chicken_rice[23][28] = 16'b10111_110111_11111;
        chicken_rice[23][29] = 16'b10111_110111_11111;
        chicken_rice[23][30] = 16'b10111_110111_11111;
        chicken_rice[23][31] = 16'b10111_110111_11111;
        chicken_rice[24][0] = 16'b10111_110111_11111;
        chicken_rice[24][1] = 16'b10111_110111_11111;
        chicken_rice[24][2] = 16'b10111_110111_11111;
        chicken_rice[24][3] = 16'b10111_110111_11111;
        chicken_rice[24][4] = 16'b10111_110111_11111;
        chicken_rice[24][5] = 16'b10111_110111_11111;
        chicken_rice[24][6] = 16'b10111_110111_11111;
        chicken_rice[24][7] = 16'b10111_110111_11111;
        chicken_rice[24][8] = 16'b10111_110111_11111;
        chicken_rice[24][9] = 16'b10111_110111_11111;
        chicken_rice[24][10] = 16'b11011_101110_01111;
        chicken_rice[24][11] = 16'b11100_110001_10001;
        chicken_rice[24][12] = 16'b11100_110001_10001;
        chicken_rice[24][13] = 16'b11011_110000_10000;
        chicken_rice[24][14] = 16'b11011_101110_01111;
        chicken_rice[24][15] = 16'b11011_101111_01111;
        chicken_rice[24][16] = 16'b11010_101101_01111;
        chicken_rice[24][17] = 16'b01110_011101_00111;
        chicken_rice[24][18] = 16'b10000_100001_01000;
        chicken_rice[24][19] = 16'b10000_100000_01000;
        chicken_rice[24][20] = 16'b10010_100101_01010;
        chicken_rice[24][21] = 16'b10001_100010_01001;
        chicken_rice[24][22] = 16'b10000_100001_01000;
        chicken_rice[24][23] = 16'b10010_100011_01001;
        chicken_rice[24][24] = 16'b01101_011011_00110;
        chicken_rice[24][25] = 16'b10111_110111_11111;
        chicken_rice[24][26] = 16'b10111_110111_11111;
        chicken_rice[24][27] = 16'b10111_110111_11111;
        chicken_rice[24][28] = 16'b10111_110111_11111;
        chicken_rice[24][29] = 16'b10111_110111_11111;
        chicken_rice[24][30] = 16'b10111_110111_11111;
        chicken_rice[24][31] = 16'b10111_110111_11111;
        chicken_rice[25][0] = 16'b10111_110111_11111;
        chicken_rice[25][1] = 16'b10111_110111_11111;
        chicken_rice[25][2] = 16'b10111_110111_11111;
        chicken_rice[25][3] = 16'b10111_110111_11111;
        chicken_rice[25][4] = 16'b10111_110111_11111;
        chicken_rice[25][5] = 16'b10111_110111_11111;
        chicken_rice[25][6] = 16'b10111_110111_11111;
        chicken_rice[25][7] = 16'b10111_110111_11111;
        chicken_rice[25][8] = 16'b10111_110111_11111;
        chicken_rice[25][9] = 16'b10111_110111_11111;
        chicken_rice[25][10] = 16'b10111_110111_11111;
        chicken_rice[25][11] = 16'b10111_110111_11111;
        chicken_rice[25][12] = 16'b10111_110111_11111;
        chicken_rice[25][13] = 16'b10111_110111_11111;
        chicken_rice[25][14] = 16'b10111_110111_11111;
        chicken_rice[25][15] = 16'b10111_110111_11111;
        chicken_rice[25][16] = 16'b10111_110111_11111;
        chicken_rice[25][17] = 16'b10111_110111_11111;
        chicken_rice[25][18] = 16'b01100_011001_00101;
        chicken_rice[25][19] = 16'b10000_100000_00111;
        chicken_rice[25][20] = 16'b10010_100100_01001;
        chicken_rice[25][21] = 16'b10101_101000_01100;
        chicken_rice[25][22] = 16'b01100_011010_00101;
        chicken_rice[25][23] = 16'b01111_011111_00111;
        chicken_rice[25][24] = 16'b10111_110111_11111;
        chicken_rice[25][25] = 16'b10111_110111_11111;
        chicken_rice[25][26] = 16'b10111_110111_11111;
        chicken_rice[25][27] = 16'b10111_110111_11111;
        chicken_rice[25][28] = 16'b10111_110111_11111;
        chicken_rice[25][29] = 16'b10111_110111_11111;
        chicken_rice[25][30] = 16'b10111_110111_11111;
        chicken_rice[25][31] = 16'b10111_110111_11111;
        chicken_rice[26][0] = 16'b10111_110111_11111;
        chicken_rice[26][1] = 16'b10111_110111_11111;
        chicken_rice[26][2] = 16'b10111_110111_11111;
        chicken_rice[26][3] = 16'b10111_110111_11111;
        chicken_rice[26][4] = 16'b10111_110111_11111;
        chicken_rice[26][5] = 16'b10111_110111_11111;
        chicken_rice[26][6] = 16'b10111_110111_11111;
        chicken_rice[26][7] = 16'b10111_110111_11111;
        chicken_rice[26][8] = 16'b10111_110111_11111;
        chicken_rice[26][9] = 16'b10111_110111_11111;
        chicken_rice[26][10] = 16'b10111_110111_11111;
        chicken_rice[26][11] = 16'b10111_110111_11111;
        chicken_rice[26][12] = 16'b10111_110111_11111;
        chicken_rice[26][13] = 16'b10111_110111_11111;
        chicken_rice[26][14] = 16'b10111_110111_11111;
        chicken_rice[26][15] = 16'b10111_110111_11111;
        chicken_rice[26][16] = 16'b10111_110111_11111;
        chicken_rice[26][17] = 16'b10111_110111_11111;
        chicken_rice[26][18] = 16'b10111_110111_11111;
        chicken_rice[26][19] = 16'b01100_011001_00101;
        chicken_rice[26][20] = 16'b01100_011010_00101;
        chicken_rice[26][21] = 16'b01101_011011_00110;
        chicken_rice[26][22] = 16'b01011_010111_00100;
        chicken_rice[26][23] = 16'b10111_110111_11111;
        chicken_rice[26][24] = 16'b10111_110111_11111;
        chicken_rice[26][25] = 16'b10111_110111_11111;
        chicken_rice[26][26] = 16'b10111_110111_11111;
        chicken_rice[26][27] = 16'b10111_110111_11111;
        chicken_rice[26][28] = 16'b10111_110111_11111;
        chicken_rice[26][29] = 16'b10111_110111_11111;
        chicken_rice[26][30] = 16'b10111_110111_11111;
        chicken_rice[26][31] = 16'b10111_110111_11111;
        chicken_rice[27][0] = 16'b10111_110111_11111;
        chicken_rice[27][1] = 16'b10111_110111_11111;
        chicken_rice[27][2] = 16'b10111_110111_11111;
        chicken_rice[27][3] = 16'b10111_110111_11111;
        chicken_rice[27][4] = 16'b10111_110111_11111;
        chicken_rice[27][5] = 16'b10111_110111_11111;
        chicken_rice[27][6] = 16'b10111_110111_11111;
        chicken_rice[27][7] = 16'b10111_110111_11111;
        chicken_rice[27][8] = 16'b10111_110111_11111;
        chicken_rice[27][9] = 16'b10111_110111_11111;
        chicken_rice[27][10] = 16'b10111_110111_11111;
        chicken_rice[27][11] = 16'b10111_110111_11111;
        chicken_rice[27][12] = 16'b10111_110111_11111;
        chicken_rice[27][13] = 16'b10111_110111_11111;
        chicken_rice[27][14] = 16'b10111_110111_11111;
        chicken_rice[27][15] = 16'b10111_110111_11111;
        chicken_rice[27][16] = 16'b10111_110111_11111;
        chicken_rice[27][17] = 16'b10111_110111_11111;
        chicken_rice[27][18] = 16'b10111_110111_11111;
        chicken_rice[27][19] = 16'b10111_110111_11111;
        chicken_rice[27][20] = 16'b10111_110111_11111;
        chicken_rice[27][21] = 16'b10111_110111_11111;
        chicken_rice[27][22] = 16'b10111_110111_11111;
        chicken_rice[27][23] = 16'b10111_110111_11111;
        chicken_rice[27][24] = 16'b10111_110111_11111;
        chicken_rice[27][25] = 16'b10111_110111_11111;
        chicken_rice[27][26] = 16'b10111_110111_11111;
        chicken_rice[27][27] = 16'b10111_110111_11111;
        chicken_rice[27][28] = 16'b10111_110111_11111;
        chicken_rice[27][29] = 16'b10111_110111_11111;
        chicken_rice[27][30] = 16'b10111_110111_11111;
        chicken_rice[27][31] = 16'b10111_110111_11111;
        chicken_rice[28][0] = 16'b10111_110111_11111;
        chicken_rice[28][1] = 16'b10111_110111_11111;
        chicken_rice[28][2] = 16'b10111_110111_11111;
        chicken_rice[28][3] = 16'b10111_110111_11111;
        chicken_rice[28][4] = 16'b10111_110111_11111;
        chicken_rice[28][5] = 16'b10111_110111_11111;
        chicken_rice[28][6] = 16'b10111_110111_11111;
        chicken_rice[28][7] = 16'b10111_110111_11111;
        chicken_rice[28][8] = 16'b10111_110111_11111;
        chicken_rice[28][9] = 16'b10111_110111_11111;
        chicken_rice[28][10] = 16'b10111_110111_11111;
        chicken_rice[28][11] = 16'b10111_110111_11111;
        chicken_rice[28][12] = 16'b10111_110111_11111;
        chicken_rice[28][13] = 16'b10111_110111_11111;
        chicken_rice[28][14] = 16'b10111_110111_11111;
        chicken_rice[28][15] = 16'b10111_110111_11111;
        chicken_rice[28][16] = 16'b10111_110111_11111;
        chicken_rice[28][17] = 16'b10111_110111_11111;
        chicken_rice[28][18] = 16'b10111_110111_11111;
        chicken_rice[28][19] = 16'b10111_110111_11111;
        chicken_rice[28][20] = 16'b10111_110111_11111;
        chicken_rice[28][21] = 16'b10111_110111_11111;
        chicken_rice[28][22] = 16'b10111_110111_11111;
        chicken_rice[28][23] = 16'b10111_110111_11111;
        chicken_rice[28][24] = 16'b10111_110111_11111;
        chicken_rice[28][25] = 16'b10111_110111_11111;
        chicken_rice[28][26] = 16'b10111_110111_11111;
        chicken_rice[28][27] = 16'b10111_110111_11111;
        chicken_rice[28][28] = 16'b10111_110111_11111;
        chicken_rice[28][29] = 16'b10111_110111_11111;
        chicken_rice[28][30] = 16'b10111_110111_11111;
        chicken_rice[28][31] = 16'b10111_110111_11111;
        chicken_rice[29][0] = 16'b10111_110111_11111;
        chicken_rice[29][1] = 16'b10111_110111_11111;
        chicken_rice[29][2] = 16'b10111_110111_11111;
        chicken_rice[29][3] = 16'b10111_110111_11111;
        chicken_rice[29][4] = 16'b10111_110111_11111;
        chicken_rice[29][5] = 16'b10111_110111_11111;
        chicken_rice[29][6] = 16'b10111_110111_11111;
        chicken_rice[29][7] = 16'b10111_110111_11111;
        chicken_rice[29][8] = 16'b10111_110111_11111;
        chicken_rice[29][9] = 16'b10111_110111_11111;
        chicken_rice[29][10] = 16'b10111_110111_11111;
        chicken_rice[29][11] = 16'b10111_110111_11111;
        chicken_rice[29][12] = 16'b10111_110111_11111;
        chicken_rice[29][13] = 16'b10111_110111_11111;
        chicken_rice[29][14] = 16'b10111_110111_11111;
        chicken_rice[29][15] = 16'b10111_110111_11111;
        chicken_rice[29][16] = 16'b10111_110111_11111;
        chicken_rice[29][17] = 16'b10111_110111_11111;
        chicken_rice[29][18] = 16'b10111_110111_11111;
        chicken_rice[29][19] = 16'b10111_110111_11111;
        chicken_rice[29][20] = 16'b10111_110111_11111;
        chicken_rice[29][21] = 16'b10111_110111_11111;
        chicken_rice[29][22] = 16'b10111_110111_11111;
        chicken_rice[29][23] = 16'b10111_110111_11111;
        chicken_rice[29][24] = 16'b10111_110111_11111;
        chicken_rice[29][25] = 16'b10111_110111_11111;
        chicken_rice[29][26] = 16'b10111_110111_11111;
        chicken_rice[29][27] = 16'b10111_110111_11111;
        chicken_rice[29][28] = 16'b10111_110111_11111;
        chicken_rice[29][29] = 16'b10111_110111_11111;
        chicken_rice[29][30] = 16'b10111_110111_11111;
        chicken_rice[29][31] = 16'b10111_110111_11111;
        chicken_rice[30][0] = 16'b10111_110111_11111;
        chicken_rice[30][1] = 16'b10111_110111_11111;
        chicken_rice[30][2] = 16'b10111_110111_11111;
        chicken_rice[30][3] = 16'b10111_110111_11111;
        chicken_rice[30][4] = 16'b10111_110111_11111;
        chicken_rice[30][5] = 16'b10111_110111_11111;
        chicken_rice[30][6] = 16'b10111_110111_11111;
        chicken_rice[30][7] = 16'b10111_110111_11111;
        chicken_rice[30][8] = 16'b10111_110111_11111;
        chicken_rice[30][9] = 16'b10111_110111_11111;
        chicken_rice[30][10] = 16'b10111_110111_11111;
        chicken_rice[30][11] = 16'b10111_110111_11111;
        chicken_rice[30][12] = 16'b10111_110111_11111;
        chicken_rice[30][13] = 16'b10111_110111_11111;
        chicken_rice[30][14] = 16'b10111_110111_11111;
        chicken_rice[30][15] = 16'b10111_110111_11111;
        chicken_rice[30][16] = 16'b10111_110111_11111;
        chicken_rice[30][17] = 16'b10111_110111_11111;
        chicken_rice[30][18] = 16'b10111_110111_11111;
        chicken_rice[30][19] = 16'b10111_110111_11111;
        chicken_rice[30][20] = 16'b10111_110111_11111;
        chicken_rice[30][21] = 16'b10111_110111_11111;
        chicken_rice[30][22] = 16'b10111_110111_11111;
        chicken_rice[30][23] = 16'b10111_110111_11111;
        chicken_rice[30][24] = 16'b10111_110111_11111;
        chicken_rice[30][25] = 16'b10111_110111_11111;
        chicken_rice[30][26] = 16'b10111_110111_11111;
        chicken_rice[30][27] = 16'b10111_110111_11111;
        chicken_rice[30][28] = 16'b10111_110111_11111;
        chicken_rice[30][29] = 16'b10111_110111_11111;
        chicken_rice[30][30] = 16'b10111_110111_11111;
        chicken_rice[30][31] = 16'b10111_110111_11111;
        chicken_rice[31][0] = 16'b10111_110111_11111;
        chicken_rice[31][1] = 16'b10111_110111_11111;
        chicken_rice[31][2] = 16'b10111_110111_11111;
        chicken_rice[31][3] = 16'b10111_110111_11111;
        chicken_rice[31][4] = 16'b10111_110111_11111;
        chicken_rice[31][5] = 16'b10111_110111_11111;
        chicken_rice[31][6] = 16'b10111_110111_11111;
        chicken_rice[31][7] = 16'b10111_110111_11111;
        chicken_rice[31][8] = 16'b10111_110111_11111;
        chicken_rice[31][9] = 16'b10111_110111_11111;
        chicken_rice[31][10] = 16'b10111_110111_11111;
        chicken_rice[31][11] = 16'b10111_110111_11111;
        chicken_rice[31][12] = 16'b10111_110111_11111;
        chicken_rice[31][13] = 16'b10111_110111_11111;
        chicken_rice[31][14] = 16'b10111_110111_11111;
        chicken_rice[31][15] = 16'b10111_110111_11111;
        chicken_rice[31][16] = 16'b10111_110111_11111;
        chicken_rice[31][17] = 16'b10111_110111_11111;
        chicken_rice[31][18] = 16'b10111_110111_11111;
        chicken_rice[31][19] = 16'b10111_110111_11111;
        chicken_rice[31][20] = 16'b10111_110111_11111;
        chicken_rice[31][21] = 16'b10111_110111_11111;
        chicken_rice[31][22] = 16'b10111_110111_11111;
        chicken_rice[31][23] = 16'b10111_110111_11111;
        chicken_rice[31][24] = 16'b10111_110111_11111;
        chicken_rice[31][25] = 16'b10111_110111_11111;
        chicken_rice[31][26] = 16'b10111_110111_11111;
        chicken_rice[31][27] = 16'b10111_110111_11111;
        chicken_rice[31][28] = 16'b10111_110111_11111;
        chicken_rice[31][29] = 16'b10111_110111_11111;
        chicken_rice[31][30] = 16'b10111_110111_11111;
        chicken_rice[31][31] = 16'b10111_110111_11111;


        
        onion_soup[0][0] = 16'b11111_101011_10101;
        onion_soup[0][1] = 16'b11111_101011_10101;
        onion_soup[0][2] = 16'b11111_101011_10101;
        onion_soup[0][3] = 16'b11111_101011_10101;
        onion_soup[0][4] = 16'b11111_101011_10101;
        onion_soup[0][5] = 16'b11111_101011_10101;
        onion_soup[0][6] = 16'b11111_101011_10101;
        onion_soup[0][7] = 16'b11111_101011_10101;
        onion_soup[0][8] = 16'b11111_101011_10101;
        onion_soup[0][9] = 16'b11111_101011_10101;
        onion_soup[0][10] = 16'b11111_101011_10101;
        onion_soup[0][11] = 16'b11111_101011_10101;
        onion_soup[0][12] = 16'b11111_101011_10101;
        onion_soup[0][13] = 16'b11111_101011_10101;
        onion_soup[0][14] = 16'b11111_101011_10101;
        onion_soup[0][15] = 16'b11111_101011_10101;
        onion_soup[0][16] = 16'b11111_101011_10101;
        onion_soup[0][17] = 16'b11111_101011_10101;
        onion_soup[0][18] = 16'b11111_101011_10101;
        onion_soup[0][19] = 16'b11111_101011_10101;
        onion_soup[0][20] = 16'b11111_101011_10101;
        onion_soup[0][21] = 16'b11111_101011_10101;
        onion_soup[0][22] = 16'b11111_101011_10101;
        onion_soup[0][23] = 16'b11111_101011_10101;
        onion_soup[0][24] = 16'b11111_101011_10101;
        onion_soup[0][25] = 16'b11111_101011_10101;
        onion_soup[0][26] = 16'b11111_101011_10101;
        onion_soup[0][27] = 16'b11111_101011_10101;
        onion_soup[0][28] = 16'b11111_101011_10101;
        onion_soup[0][29] = 16'b11111_101011_10101;
        onion_soup[0][30] = 16'b11111_101011_10101;
        onion_soup[0][31] = 16'b11111_101011_10101;
        onion_soup[1][0] = 16'b11111_101011_10101;
        onion_soup[1][1] = 16'b11111_101011_10101;
        onion_soup[1][2] = 16'b11111_101011_10101;
        onion_soup[1][3] = 16'b11111_101011_10101;
        onion_soup[1][4] = 16'b11111_101011_10101;
        onion_soup[1][5] = 16'b11111_101011_10101;
        onion_soup[1][6] = 16'b11111_101011_10101;
        onion_soup[1][7] = 16'b11111_101011_10101;
        onion_soup[1][8] = 16'b11111_101011_10101;
        onion_soup[1][9] = 16'b11111_101011_10101;
        onion_soup[1][10] = 16'b11111_101011_10101;
        onion_soup[1][11] = 16'b11111_101011_10101;
        onion_soup[1][12] = 16'b11111_101011_10101;
        onion_soup[1][13] = 16'b11111_101011_10101;
        onion_soup[1][14] = 16'b11111_101011_10101;
        onion_soup[1][15] = 16'b11111_101011_10101;
        onion_soup[1][16] = 16'b11111_101011_10101;
        onion_soup[1][17] = 16'b11111_101011_10101;
        onion_soup[1][18] = 16'b11111_101011_10101;
        onion_soup[1][19] = 16'b11111_101011_10101;
        onion_soup[1][20] = 16'b11111_101011_10101;
        onion_soup[1][21] = 16'b11111_101011_10101;
        onion_soup[1][22] = 16'b11111_101011_10101;
        onion_soup[1][23] = 16'b11111_101011_10101;
        onion_soup[1][24] = 16'b11111_101011_10101;
        onion_soup[1][25] = 16'b11111_101011_10101;
        onion_soup[1][26] = 16'b11111_101011_10101;
        onion_soup[1][27] = 16'b11111_101011_10101;
        onion_soup[1][28] = 16'b11111_101011_10101;
        onion_soup[1][29] = 16'b11111_101011_10101;
        onion_soup[1][30] = 16'b11111_101011_10101;
        onion_soup[1][31] = 16'b11111_101011_10101;
        onion_soup[2][0] = 16'b11111_101011_10101;
        onion_soup[2][1] = 16'b11111_101011_10101;
        onion_soup[2][2] = 16'b11111_101011_10101;
        onion_soup[2][3] = 16'b11111_101011_10101;
        onion_soup[2][4] = 16'b11111_101011_10101;
        onion_soup[2][5] = 16'b11111_101011_10101;
        onion_soup[2][6] = 16'b11111_101011_10101;
        onion_soup[2][7] = 16'b11111_101011_10101;
        onion_soup[2][8] = 16'b11111_101011_10101;
        onion_soup[2][9] = 16'b11111_101011_10101;
        onion_soup[2][10] = 16'b11111_101011_10101;
        onion_soup[2][11] = 16'b11111_101011_10101;
        onion_soup[2][12] = 16'b11111_101011_10101;
        onion_soup[2][13] = 16'b11111_101011_10101;
        onion_soup[2][14] = 16'b11111_101011_10101;
        onion_soup[2][15] = 16'b11111_101011_10101;
        onion_soup[2][16] = 16'b11111_101011_10101;
        onion_soup[2][17] = 16'b11111_101011_10101;
        onion_soup[2][18] = 16'b11111_101011_10101;
        onion_soup[2][19] = 16'b11111_101011_10101;
        onion_soup[2][20] = 16'b11111_101011_10101;
        onion_soup[2][21] = 16'b11111_101011_10101;
        onion_soup[2][22] = 16'b11111_101011_10101;
        onion_soup[2][23] = 16'b11111_101011_10101;
        onion_soup[2][24] = 16'b11111_101011_10101;
        onion_soup[2][25] = 16'b11111_101011_10101;
        onion_soup[2][26] = 16'b11111_101011_10101;
        onion_soup[2][27] = 16'b11111_101011_10101;
        onion_soup[2][28] = 16'b11111_101011_10101;
        onion_soup[2][29] = 16'b11111_101011_10101;
        onion_soup[2][30] = 16'b11111_101011_10101;
        onion_soup[2][31] = 16'b11111_101011_10101;
        onion_soup[3][0] = 16'b11111_101011_10101;
        onion_soup[3][1] = 16'b11111_101011_10101;
        onion_soup[3][2] = 16'b11111_101011_10101;
        onion_soup[3][3] = 16'b11111_101011_10101;
        onion_soup[3][4] = 16'b11111_101011_10101;
        onion_soup[3][5] = 16'b11111_101011_10101;
        onion_soup[3][6] = 16'b11111_101011_10101;
        onion_soup[3][7] = 16'b11111_101011_10101;
        onion_soup[3][8] = 16'b11111_101011_10101;
        onion_soup[3][9] = 16'b11111_101011_10101;
        onion_soup[3][10] = 16'b11111_101011_10101;
        onion_soup[3][11] = 16'b11111_101011_10101;
        onion_soup[3][12] = 16'b11111_101011_10101;
        onion_soup[3][13] = 16'b11111_101011_10101;
        onion_soup[3][14] = 16'b11111_101011_10101;
        onion_soup[3][15] = 16'b11111_101011_10101;
        onion_soup[3][16] = 16'b11111_101011_10101;
        onion_soup[3][17] = 16'b11111_101011_10101;
        onion_soup[3][18] = 16'b11111_101011_10101;
        onion_soup[3][19] = 16'b11111_101011_10101;
        onion_soup[3][20] = 16'b11111_101011_10101;
        onion_soup[3][21] = 16'b11111_101011_10101;
        onion_soup[3][22] = 16'b11111_101011_10101;
        onion_soup[3][23] = 16'b11111_101011_10101;
        onion_soup[3][24] = 16'b11111_101011_10101;
        onion_soup[3][25] = 16'b11111_101011_10101;
        onion_soup[3][26] = 16'b11111_101011_10101;
        onion_soup[3][27] = 16'b11111_101011_10101;
        onion_soup[3][28] = 16'b11111_101011_10101;
        onion_soup[3][29] = 16'b11111_101011_10101;
        onion_soup[3][30] = 16'b11111_101011_10101;
        onion_soup[3][31] = 16'b11111_101011_10101;
        onion_soup[4][0] = 16'b11111_101011_10101;
        onion_soup[4][1] = 16'b11111_101011_10101;
        onion_soup[4][2] = 16'b11111_101011_10101;
        onion_soup[4][3] = 16'b11111_101011_10101;
        onion_soup[4][4] = 16'b11111_101011_10101;
        onion_soup[4][5] = 16'b11111_101011_10101;
        onion_soup[4][6] = 16'b11111_101011_10101;
        onion_soup[4][7] = 16'b11111_101011_10101;
        onion_soup[4][8] = 16'b11111_101011_10101;
        onion_soup[4][9] = 16'b11111_101011_10101;
        onion_soup[4][10] = 16'b11111_101011_10101;
        onion_soup[4][11] = 16'b11111_101011_10101;
        onion_soup[4][12] = 16'b11111_101011_10101;
        onion_soup[4][13] = 16'b11111_101011_10101;
        onion_soup[4][14] = 16'b11111_101011_10101;
        onion_soup[4][15] = 16'b11111_101011_10101;
        onion_soup[4][16] = 16'b11111_101011_10101;
        onion_soup[4][17] = 16'b11111_101011_10101;
        onion_soup[4][18] = 16'b11111_101011_10101;
        onion_soup[4][19] = 16'b11111_101011_10101;
        onion_soup[4][20] = 16'b11111_101011_10101;
        onion_soup[4][21] = 16'b11111_101011_10101;
        onion_soup[4][22] = 16'b11111_101011_10101;
        onion_soup[4][23] = 16'b11111_101011_10101;
        onion_soup[4][24] = 16'b11111_101011_10101;
        onion_soup[4][25] = 16'b11111_101011_10101;
        onion_soup[4][26] = 16'b11111_101011_10101;
        onion_soup[4][27] = 16'b11111_101011_10101;
        onion_soup[4][28] = 16'b11111_101011_10101;
        onion_soup[4][29] = 16'b11111_101011_10101;
        onion_soup[4][30] = 16'b11111_101011_10101;
        onion_soup[4][31] = 16'b11111_101011_10101;
        onion_soup[5][0] = 16'b11111_101011_10101;
        onion_soup[5][1] = 16'b11111_101011_10101;
        onion_soup[5][2] = 16'b11111_101011_10101;
        onion_soup[5][3] = 16'b11111_101011_10101;
        onion_soup[5][4] = 16'b11111_101011_10101;
        onion_soup[5][5] = 16'b11111_101011_10101;
        onion_soup[5][6] = 16'b11111_101011_10101;
        onion_soup[5][7] = 16'b11111_101011_10101;
        onion_soup[5][8] = 16'b11111_101011_10101;
        onion_soup[5][9] = 16'b11111_101011_10101;
        onion_soup[5][10] = 16'b11111_101011_10101;
        onion_soup[5][11] = 16'b11111_101011_10101;
        onion_soup[5][12] = 16'b11111_101011_10101;
        onion_soup[5][13] = 16'b11111_101011_10101;
        onion_soup[5][14] = 16'b11111_101011_10101;
        onion_soup[5][15] = 16'b11111_101011_10101;
        onion_soup[5][16] = 16'b11111_101011_10101;
        onion_soup[5][17] = 16'b11111_101011_10101;
        onion_soup[5][18] = 16'b11111_101011_10101;
        onion_soup[5][19] = 16'b11111_101011_10101;
        onion_soup[5][20] = 16'b11111_101011_10101;
        onion_soup[5][21] = 16'b11111_101011_10101;
        onion_soup[5][22] = 16'b11111_101011_10101;
        onion_soup[5][23] = 16'b11111_101011_10101;
        onion_soup[5][24] = 16'b11111_101011_10101;
        onion_soup[5][25] = 16'b11111_101011_10101;
        onion_soup[5][26] = 16'b11111_101011_10101;
        onion_soup[5][27] = 16'b11111_101011_10101;
        onion_soup[5][28] = 16'b11111_101011_10101;
        onion_soup[5][29] = 16'b11111_101011_10101;
        onion_soup[5][30] = 16'b11111_101011_10101;
        onion_soup[5][31] = 16'b11111_101011_10101;
        onion_soup[6][0] = 16'b11111_101011_10101;
        onion_soup[6][1] = 16'b11111_101011_10101;
        onion_soup[6][2] = 16'b11111_101011_10101;
        onion_soup[6][3] = 16'b11111_101011_10101;
        onion_soup[6][4] = 16'b11111_101011_10101;
        onion_soup[6][5] = 16'b11111_101011_10101;
        onion_soup[6][6] = 16'b11111_101011_10101;
        onion_soup[6][7] = 16'b11111_101011_10101;
        onion_soup[6][8] = 16'b11111_101011_10101;
        onion_soup[6][9] = 16'b11111_101011_10101;
        onion_soup[6][10] = 16'b11111_101011_10101;
        onion_soup[6][11] = 16'b11111_101011_10101;
        onion_soup[6][12] = 16'b10001_010100_00011;
        onion_soup[6][13] = 16'b10001_010101_00011;
        onion_soup[6][14] = 16'b10101_011011_00100;
        onion_soup[6][15] = 16'b10010_010110_00011;
        onion_soup[6][16] = 16'b10010_010101_00011;
        onion_soup[6][17] = 16'b10000_010100_00010;
        onion_soup[6][18] = 16'b10010_010110_00011;
        onion_soup[6][19] = 16'b10011_011000_00100;
        onion_soup[6][20] = 16'b10001_010100_00010;
        onion_soup[6][21] = 16'b11111_101011_10101;
        onion_soup[6][22] = 16'b11111_101011_10101;
        onion_soup[6][23] = 16'b11111_101011_10101;
        onion_soup[6][24] = 16'b11111_101011_10101;
        onion_soup[6][25] = 16'b11111_101011_10101;
        onion_soup[6][26] = 16'b11111_101011_10101;
        onion_soup[6][27] = 16'b11111_101011_10101;
        onion_soup[6][28] = 16'b11111_101011_10101;
        onion_soup[6][29] = 16'b11111_101011_10101;
        onion_soup[6][30] = 16'b11111_101011_10101;
        onion_soup[6][31] = 16'b11111_101011_10101;
        onion_soup[7][0] = 16'b11111_101011_10101;
        onion_soup[7][1] = 16'b11111_101011_10101;
        onion_soup[7][2] = 16'b11111_101011_10101;
        onion_soup[7][3] = 16'b11111_101011_10101;
        onion_soup[7][4] = 16'b11111_101011_10101;
        onion_soup[7][5] = 16'b11111_101011_10101;
        onion_soup[7][6] = 16'b11111_101011_10101;
        onion_soup[7][7] = 16'b11111_101011_10101;
        onion_soup[7][8] = 16'b11111_101011_10101;
        onion_soup[7][9] = 16'b11111_101011_10101;
        onion_soup[7][10] = 16'b10000_010011_00010;
        onion_soup[7][11] = 16'b01111_010010_00010;
        onion_soup[7][12] = 16'b10011_011010_00101;
        onion_soup[7][13] = 16'b10001_010110_00011;
        onion_soup[7][14] = 16'b10111_011111_00110;
        onion_soup[7][15] = 16'b10010_010110_00011;
        onion_soup[7][16] = 16'b10110_011101_00110;
        onion_soup[7][17] = 16'b11000_100011_01000;
        onion_soup[7][18] = 16'b01111_010010_00010;
        onion_soup[7][19] = 16'b10011_011001_00100;
        onion_soup[7][20] = 16'b01111_010010_00010;
        onion_soup[7][21] = 16'b10000_010011_00010;
        onion_soup[7][22] = 16'b10000_010011_00011;
        onion_soup[7][23] = 16'b11111_101011_10101;
        onion_soup[7][24] = 16'b11111_101011_10101;
        onion_soup[7][25] = 16'b11111_101011_10101;
        onion_soup[7][26] = 16'b11111_101011_10101;
        onion_soup[7][27] = 16'b11111_101011_10101;
        onion_soup[7][28] = 16'b11111_101011_10101;
        onion_soup[7][29] = 16'b11111_101011_10101;
        onion_soup[7][30] = 16'b11111_101011_10101;
        onion_soup[7][31] = 16'b11111_101011_10101;
        onion_soup[8][0] = 16'b11111_101011_10101;
        onion_soup[8][1] = 16'b11111_101011_10101;
        onion_soup[8][2] = 16'b11111_101011_10101;
        onion_soup[8][3] = 16'b11111_101011_10101;
        onion_soup[8][4] = 16'b11111_101011_10101;
        onion_soup[8][5] = 16'b11111_101011_10101;
        onion_soup[8][6] = 16'b11111_101011_10101;
        onion_soup[8][7] = 16'b11111_101011_10101;
        onion_soup[8][8] = 16'b10100_011001_00100;
        onion_soup[8][9] = 16'b10011_011001_00100;
        onion_soup[8][10] = 16'b10111_100000_00111;
        onion_soup[8][11] = 16'b10100_011010_00101;
        onion_soup[8][12] = 16'b10100_011010_00101;
        onion_soup[8][13] = 16'b10011_011000_00100;
        onion_soup[8][14] = 16'b10011_011000_00100;
        onion_soup[8][15] = 16'b11010_100110_01001;
        onion_soup[8][16] = 16'b10100_011010_00101;
        onion_soup[8][17] = 16'b10110_011101_00101;
        onion_soup[8][18] = 16'b10011_010111_00100;
        onion_soup[8][19] = 16'b10111_011111_00110;
        onion_soup[8][20] = 16'b10000_010011_00011;
        onion_soup[8][21] = 16'b10100_011010_00100;
        onion_soup[8][22] = 16'b10100_011010_00100;
        onion_soup[8][23] = 16'b10000_010011_00010;
        onion_soup[8][24] = 16'b11111_101011_10101;
        onion_soup[8][25] = 16'b11111_101011_10101;
        onion_soup[8][26] = 16'b11111_101011_10101;
        onion_soup[8][27] = 16'b11111_101011_10101;
        onion_soup[8][28] = 16'b11111_101011_10101;
        onion_soup[8][29] = 16'b11111_101011_10101;
        onion_soup[8][30] = 16'b11111_101011_10101;
        onion_soup[8][31] = 16'b11111_101011_10101;
        onion_soup[9][0] = 16'b11111_101011_10101;
        onion_soup[9][1] = 16'b11111_101011_10101;
        onion_soup[9][2] = 16'b11111_101011_10101;
        onion_soup[9][3] = 16'b11111_101011_10101;
        onion_soup[9][4] = 16'b11111_101011_10101;
        onion_soup[9][5] = 16'b11111_101011_10101;
        onion_soup[9][6] = 16'b11111_101011_10101;
        onion_soup[9][7] = 16'b10001_010100_00011;
        onion_soup[9][8] = 16'b10100_011011_00101;
        onion_soup[9][9] = 16'b11001_100100_01001;
        onion_soup[9][10] = 16'b11001_100101_01001;
        onion_soup[9][11] = 16'b10101_011101_00110;
        onion_soup[9][12] = 16'b10110_011101_00110;
        onion_soup[9][13] = 16'b10100_011011_00101;
        onion_soup[9][14] = 16'b11010_100110_01001;
        onion_soup[9][15] = 16'b10100_011010_00101;
        onion_soup[9][16] = 16'b10010_010110_00011;
        onion_soup[9][17] = 16'b10111_011111_00110;
        onion_soup[9][18] = 16'b10110_011101_00101;
        onion_soup[9][19] = 16'b10101_011101_00110;
        onion_soup[9][20] = 16'b01110_001111_00010;
        onion_soup[9][21] = 16'b10101_011011_00101;
        onion_soup[9][22] = 16'b10110_011101_00110;
        onion_soup[9][23] = 16'b10100_011001_00101;
        onion_soup[9][24] = 16'b10011_011000_00100;
        onion_soup[9][25] = 16'b11111_101011_10101;
        onion_soup[9][26] = 16'b11111_101011_10101;
        onion_soup[9][27] = 16'b11111_101011_10101;
        onion_soup[9][28] = 16'b11111_101011_10101;
        onion_soup[9][29] = 16'b11111_101011_10101;
        onion_soup[9][30] = 16'b11111_101011_10101;
        onion_soup[9][31] = 16'b11111_101011_10101;
        onion_soup[10][0] = 16'b11111_101011_10101;
        onion_soup[10][1] = 16'b11111_101011_10101;
        onion_soup[10][2] = 16'b11111_101011_10101;
        onion_soup[10][3] = 16'b11111_101011_10101;
        onion_soup[10][4] = 16'b11111_101011_10101;
        onion_soup[10][5] = 16'b11111_101011_10101;
        onion_soup[10][6] = 16'b01100_001101_00001;
        onion_soup[10][7] = 16'b10010_010111_00100;
        onion_soup[10][8] = 16'b10101_011100_00101;
        onion_soup[10][9] = 16'b10110_011101_00110;
        onion_soup[10][10] = 16'b11011_101010_01011;
        onion_soup[10][11] = 16'b10110_011110_00110;
        onion_soup[10][12] = 16'b01100_001101_00001;
        onion_soup[10][13] = 16'b10000_010011_00010;
        onion_soup[10][14] = 16'b01011_001011_00001;
        onion_soup[10][15] = 16'b01110_010000_00010;
        onion_soup[10][16] = 16'b01100_001101_00001;
        onion_soup[10][17] = 16'b10010_010111_00011;
        onion_soup[10][18] = 16'b01110_010000_00001;
        onion_soup[10][19] = 16'b10000_010011_00010;
        onion_soup[10][20] = 16'b10000_010011_00010;
        onion_soup[10][21] = 16'b01111_010010_00010;
        onion_soup[10][22] = 16'b10101_011100_00101;
        onion_soup[10][23] = 16'b10111_100000_00111;
        onion_soup[10][24] = 16'b10001_010101_00011;
        onion_soup[10][25] = 16'b10011_010111_00011;
        onion_soup[10][26] = 16'b10001_010110_00011;
        onion_soup[10][27] = 16'b11111_101011_10101;
        onion_soup[10][28] = 16'b11111_101011_10101;
        onion_soup[10][29] = 16'b11111_101011_10101;
        onion_soup[10][30] = 16'b11111_101011_10101;
        onion_soup[10][31] = 16'b11111_101011_10101;
        onion_soup[11][0] = 16'b11111_101011_10101;
        onion_soup[11][1] = 16'b11111_101011_10101;
        onion_soup[11][2] = 16'b11111_101011_10101;
        onion_soup[11][3] = 16'b11111_101011_10101;
        onion_soup[11][4] = 16'b11111_101011_10101;
        onion_soup[11][5] = 16'b10001_010101_00011;
        onion_soup[11][6] = 16'b10100_011010_00101;
        onion_soup[11][7] = 16'b10110_011101_00110;
        onion_soup[11][8] = 16'b10100_011010_00101;
        onion_soup[11][9] = 16'b01101_001111_00001;
        onion_soup[11][10] = 16'b10010_010110_00011;
        onion_soup[11][11] = 16'b10010_010110_00011;
        onion_soup[11][12] = 16'b10000_010100_00011;
        onion_soup[11][13] = 16'b10000_010010_00010;
        onion_soup[11][14] = 16'b10011_011000_00011;
        onion_soup[11][15] = 16'b10100_011001_00011;
        onion_soup[11][16] = 16'b10010_010101_00011;
        onion_soup[11][17] = 16'b10001_010101_00011;
        onion_soup[11][18] = 16'b10000_010011_00010;
        onion_soup[11][19] = 16'b10000_010011_00010;
        onion_soup[11][20] = 16'b01111_010001_00010;
        onion_soup[11][21] = 16'b01110_010001_00010;
        onion_soup[11][22] = 16'b10000_010011_00010;
        onion_soup[11][23] = 16'b01101_001111_00001;
        onion_soup[11][24] = 16'b10100_011001_00100;
        onion_soup[11][25] = 16'b10011_011000_00100;
        onion_soup[11][26] = 16'b01111_010010_00011;
        onion_soup[11][27] = 16'b11111_101011_10101;
        onion_soup[11][28] = 16'b11111_101011_10101;
        onion_soup[11][29] = 16'b11111_101011_10101;
        onion_soup[11][30] = 16'b11111_101011_10101;
        onion_soup[11][31] = 16'b11111_101011_10101;
        onion_soup[12][0] = 16'b11111_101011_10101;
        onion_soup[12][1] = 16'b11111_101011_10101;
        onion_soup[12][2] = 16'b11111_101011_10101;
        onion_soup[12][3] = 16'b11111_101011_10101;
        onion_soup[12][4] = 16'b11111_101011_10101;
        onion_soup[12][5] = 16'b10011_011010_00101;
        onion_soup[12][6] = 16'b10100_011010_00100;
        onion_soup[12][7] = 16'b01101_001111_00001;
        onion_soup[12][8] = 16'b01111_010001_00010;
        onion_soup[12][9] = 16'b01100_001100_00001;
        onion_soup[12][10] = 16'b01101_001110_00001;
        onion_soup[12][11] = 16'b01111_010001_00010;
        onion_soup[12][12] = 16'b01010_001001_00000;
        onion_soup[12][13] = 16'b01000_001000_00000;
        onion_soup[12][14] = 16'b01100_001100_00001;
        onion_soup[12][15] = 16'b01000_000111_00000;
        onion_soup[12][16] = 16'b01111_010000_00001;
        onion_soup[12][17] = 16'b00111_000111_00000;
        onion_soup[12][18] = 16'b01011_001011_00001;
        onion_soup[12][19] = 16'b01101_001101_00001;
        onion_soup[12][20] = 16'b01101_001110_00001;
        onion_soup[12][21] = 16'b10010_010101_00011;
        onion_soup[12][22] = 16'b01110_010000_00010;
        onion_soup[12][23] = 16'b10010_010111_00011;
        onion_soup[12][24] = 16'b01011_001011_00001;
        onion_soup[12][25] = 16'b10011_011001_00100;
        onion_soup[12][26] = 16'b01001_001001_00001;
        onion_soup[12][27] = 16'b11111_101011_10101;
        onion_soup[12][28] = 16'b11111_101011_10101;
        onion_soup[12][29] = 16'b11111_101011_10101;
        onion_soup[12][30] = 16'b11111_101011_10101;
        onion_soup[12][31] = 16'b11111_101011_10101;
        onion_soup[13][0] = 16'b11111_101011_10101;
        onion_soup[13][1] = 16'b11111_101011_10101;
        onion_soup[13][2] = 16'b11111_101011_10101;
        onion_soup[13][3] = 16'b11111_101011_10101;
        onion_soup[13][4] = 16'b11000_100001_00110;
        onion_soup[13][5] = 16'b01101_001111_00001;
        onion_soup[13][6] = 16'b01110_010001_00010;
        onion_soup[13][7] = 16'b10100_011010_00100;
        onion_soup[13][8] = 16'b01100_001101_00001;
        onion_soup[13][9] = 16'b01001_001001_00000;
        onion_soup[13][10] = 16'b01011_001011_00001;
        onion_soup[13][11] = 16'b01001_001000_00000;
        onion_soup[13][12] = 16'b01010_001011_00001;
        onion_soup[13][13] = 16'b10011_010111_00011;
        onion_soup[13][14] = 16'b01000_001000_00000;
        onion_soup[13][15] = 16'b01011_001011_00001;
        onion_soup[13][16] = 16'b01111_010001_00010;
        onion_soup[13][17] = 16'b01100_001110_00001;
        onion_soup[13][18] = 16'b01101_001110_00001;
        onion_soup[13][19] = 16'b01101_001110_00001;
        onion_soup[13][20] = 16'b01011_001011_00000;
        onion_soup[13][21] = 16'b01110_001111_00001;
        onion_soup[13][22] = 16'b01101_001111_00001;
        onion_soup[13][23] = 16'b01100_001101_00001;
        onion_soup[13][24] = 16'b10001_010101_00011;
        onion_soup[13][25] = 16'b10000_010011_00010;
        onion_soup[13][26] = 16'b01111_010010_00010;
        onion_soup[13][27] = 16'b10010_010111_00011;
        onion_soup[13][28] = 16'b11111_101011_10101;
        onion_soup[13][29] = 16'b11111_101011_10101;
        onion_soup[13][30] = 16'b11111_101011_10101;
        onion_soup[13][31] = 16'b11111_101011_10101;
        onion_soup[14][0] = 16'b11111_101011_10101;
        onion_soup[14][1] = 16'b11111_101011_10101;
        onion_soup[14][2] = 16'b11111_101011_10101;
        onion_soup[14][3] = 16'b11111_101011_10101;
        onion_soup[14][4] = 16'b10011_011000_00100;
        onion_soup[14][5] = 16'b01001_001001_00001;
        onion_soup[14][6] = 16'b01110_010000_00001;
        onion_soup[14][7] = 16'b01011_001100_00001;
        onion_soup[14][8] = 16'b01011_001011_00001;
        onion_soup[14][9] = 16'b01110_001111_00001;
        onion_soup[14][10] = 16'b01100_001100_00001;
        onion_soup[14][11] = 16'b01100_001101_00001;
        onion_soup[14][12] = 16'b01011_001100_00001;
        onion_soup[14][13] = 16'b01100_001100_00001;
        onion_soup[14][14] = 16'b01001_001001_00000;
        onion_soup[14][15] = 16'b01100_001101_00001;
        onion_soup[14][16] = 16'b01001_001000_00000;
        onion_soup[14][17] = 16'b10011_011010_00101;
        onion_soup[14][18] = 16'b10110_011111_00111;
        onion_soup[14][19] = 16'b01101_001110_00001;
        onion_soup[14][20] = 16'b01100_001100_00001;
        onion_soup[14][21] = 16'b01011_001100_00001;
        onion_soup[14][22] = 16'b01100_001101_00001;
        onion_soup[14][23] = 16'b01100_001100_00001;
        onion_soup[14][24] = 16'b01010_001011_00001;
        onion_soup[14][25] = 16'b01110_010000_00010;
        onion_soup[14][26] = 16'b10000_010010_00010;
        onion_soup[14][27] = 16'b10011_011001_00100;
        onion_soup[14][28] = 16'b11111_101011_10101;
        onion_soup[14][29] = 16'b11111_101011_10101;
        onion_soup[14][30] = 16'b11111_101011_10101;
        onion_soup[14][31] = 16'b11111_101011_10101;
        onion_soup[15][0] = 16'b11111_101011_10101;
        onion_soup[15][1] = 16'b11111_101011_10101;
        onion_soup[15][2] = 16'b11111_101011_10101;
        onion_soup[15][3] = 16'b11111_101011_10101;
        onion_soup[15][4] = 16'b01101_001110_00001;
        onion_soup[15][5] = 16'b01110_001111_00001;
        onion_soup[15][6] = 16'b10000_010010_00010;
        onion_soup[15][7] = 16'b01101_001110_00001;
        onion_soup[15][8] = 16'b11000_100001_00111;
        onion_soup[15][9] = 16'b11010_100111_01011;
        onion_soup[15][10] = 16'b11000_100010_00111;
        onion_soup[15][11] = 16'b01011_001011_00001;
        onion_soup[15][12] = 16'b01101_001111_00001;
        onion_soup[15][13] = 16'b01011_001100_00001;
        onion_soup[15][14] = 16'b10000_010011_00010;
        onion_soup[15][15] = 16'b01001_001000_00000;
        onion_soup[15][16] = 16'b01111_010001_00010;
        onion_soup[15][17] = 16'b10000_010010_00010;
        onion_soup[15][18] = 16'b01101_001110_00001;
        onion_soup[15][19] = 16'b01110_010000_00001;
        onion_soup[15][20] = 16'b01110_010000_00001;
        onion_soup[15][21] = 16'b01010_001010_00001;
        onion_soup[15][22] = 16'b01111_010001_00010;
        onion_soup[15][23] = 16'b01101_001111_00001;
        onion_soup[15][24] = 16'b01010_001010_00001;
        onion_soup[15][25] = 16'b01111_010000_00001;
        onion_soup[15][26] = 16'b01111_010001_00010;
        onion_soup[15][27] = 16'b10000_010011_00010;
        onion_soup[15][28] = 16'b11111_101011_10101;
        onion_soup[15][29] = 16'b11111_101011_10101;
        onion_soup[15][30] = 16'b11111_101011_10101;
        onion_soup[15][31] = 16'b11111_101011_10101;
        onion_soup[16][0] = 16'b11111_101011_10101;
        onion_soup[16][1] = 16'b11111_101011_10101;
        onion_soup[16][2] = 16'b11111_101011_10101;
        onion_soup[16][3] = 16'b11111_101011_10101;
        onion_soup[16][4] = 16'b10001_010100_00010;
        onion_soup[16][5] = 16'b10011_011000_00011;
        onion_soup[16][6] = 16'b01011_001100_00001;
        onion_soup[16][7] = 16'b01101_001101_00001;
        onion_soup[16][8] = 16'b01110_010000_00001;
        onion_soup[16][9] = 16'b01101_001110_00001;
        onion_soup[16][10] = 16'b01010_001011_00001;
        onion_soup[16][11] = 16'b01111_010001_00001;
        onion_soup[16][12] = 16'b01110_010000_00001;
        onion_soup[16][13] = 16'b01011_001100_00001;
        onion_soup[16][14] = 16'b01101_001110_00010;
        onion_soup[16][15] = 16'b10111_100000_00111;
        onion_soup[16][16] = 16'b11011_100111_01001;
        onion_soup[16][17] = 16'b10000_010010_00010;
        onion_soup[16][18] = 16'b01100_001110_00001;
        onion_soup[16][19] = 16'b01011_001011_00001;
        onion_soup[16][20] = 16'b01010_001001_00000;
        onion_soup[16][21] = 16'b10100_011001_00100;
        onion_soup[16][22] = 16'b10111_100001_01000;
        onion_soup[16][23] = 16'b11011_101101_01110;
        onion_soup[16][24] = 16'b01110_001111_00001;
        onion_soup[16][25] = 16'b01101_001101_00001;
        onion_soup[16][26] = 16'b10000_010100_00011;
        onion_soup[16][27] = 16'b01110_010000_00001;
        onion_soup[16][28] = 16'b11111_101011_10101;
        onion_soup[16][29] = 16'b11111_101011_10101;
        onion_soup[16][30] = 16'b11111_101011_10101;
        onion_soup[16][31] = 16'b11111_101011_10101;
        onion_soup[17][0] = 16'b11111_101011_10101;
        onion_soup[17][1] = 16'b11111_101011_10101;
        onion_soup[17][2] = 16'b11111_101011_10101;
        onion_soup[17][3] = 16'b11111_101011_10101;
        onion_soup[17][4] = 16'b01101_001110_00001;
        onion_soup[17][5] = 16'b10000_010100_00011;
        onion_soup[17][6] = 16'b01010_001011_00001;
        onion_soup[17][7] = 16'b01011_001011_00001;
        onion_soup[17][8] = 16'b01100_001101_00001;
        onion_soup[17][9] = 16'b01110_001111_00001;
        onion_soup[17][10] = 16'b10010_010111_00011;
        onion_soup[17][11] = 16'b10010_010110_00011;
        onion_soup[17][12] = 16'b01110_001111_00001;
        onion_soup[17][13] = 16'b01101_001110_00001;
        onion_soup[17][14] = 16'b10001_010100_00010;
        onion_soup[17][15] = 16'b01111_010001_00010;
        onion_soup[17][16] = 16'b01111_010001_00010;
        onion_soup[17][17] = 16'b10001_010100_00010;
        onion_soup[17][18] = 16'b01100_001101_00001;
        onion_soup[17][19] = 16'b10001_010101_00011;
        onion_soup[17][20] = 16'b01110_010000_00010;
        onion_soup[17][21] = 16'b01101_001110_00001;
        onion_soup[17][22] = 16'b01110_001111_00001;
        onion_soup[17][23] = 16'b01011_001011_00001;
        onion_soup[17][24] = 16'b01011_001100_00001;
        onion_soup[17][25] = 16'b01111_010001_00010;
        onion_soup[17][26] = 16'b01111_010010_00010;
        onion_soup[17][27] = 16'b10001_010110_00011;
        onion_soup[17][28] = 16'b11111_101011_10101;
        onion_soup[17][29] = 16'b11111_101011_10101;
        onion_soup[17][30] = 16'b11111_101011_10101;
        onion_soup[17][31] = 16'b11111_101011_10101;
        onion_soup[18][0] = 16'b11111_101011_10101;
        onion_soup[18][1] = 16'b11111_101011_10101;
        onion_soup[18][2] = 16'b11111_101011_10101;
        onion_soup[18][3] = 16'b11111_101011_10101;
        onion_soup[18][4] = 16'b01110_001111_00010;
        onion_soup[18][5] = 16'b10111_100001_00111;
        onion_soup[18][6] = 16'b01001_001000_00000;
        onion_soup[18][7] = 16'b01011_001100_00001;
        onion_soup[18][8] = 16'b01010_001010_00001;
        onion_soup[18][9] = 16'b01011_001011_00000;
        onion_soup[18][10] = 16'b01110_010000_00010;
        onion_soup[18][11] = 16'b11010_101001_01101;
        onion_soup[18][12] = 16'b10011_011001_00100;
        onion_soup[18][13] = 16'b01100_001101_00001;
        onion_soup[18][14] = 16'b01111_010001_00010;
        onion_soup[18][15] = 16'b10001_010101_00010;
        onion_soup[18][16] = 16'b01110_010000_00001;
        onion_soup[18][17] = 16'b01101_001111_00001;
        onion_soup[18][18] = 16'b10001_011000_00110;
        onion_soup[18][19] = 16'b10111_100000_00111;
        onion_soup[18][20] = 16'b10111_100001_01000;
        onion_soup[18][21] = 16'b01100_001101_00001;
        onion_soup[18][22] = 16'b01100_001100_00001;
        onion_soup[18][23] = 16'b01011_001011_00001;
        onion_soup[18][24] = 16'b01110_001111_00001;
        onion_soup[18][25] = 16'b10000_010100_00010;
        onion_soup[18][26] = 16'b10011_011001_00101;
        onion_soup[18][27] = 16'b10111_100000_00110;
        onion_soup[18][28] = 16'b11111_101011_10101;
        onion_soup[18][29] = 16'b11111_101011_10101;
        onion_soup[18][30] = 16'b11111_101011_10101;
        onion_soup[18][31] = 16'b11111_101011_10101;
        onion_soup[19][0] = 16'b11111_101011_10101;
        onion_soup[19][1] = 16'b11111_101011_10101;
        onion_soup[19][2] = 16'b11111_101011_10101;
        onion_soup[19][3] = 16'b11111_101011_10101;
        onion_soup[19][4] = 16'b11111_101011_10101;
        onion_soup[19][5] = 16'b01101_001111_00010;
        onion_soup[19][6] = 16'b10101_011100_00101;
        onion_soup[19][7] = 16'b01011_001011_00001;
        onion_soup[19][8] = 16'b01101_001110_00001;
        onion_soup[19][9] = 16'b01011_001011_00001;
        onion_soup[19][10] = 16'b01011_001011_00001;
        onion_soup[19][11] = 16'b01111_010001_00010;
        onion_soup[19][12] = 16'b10000_010010_00010;
        onion_soup[19][13] = 16'b01011_001100_00001;
        onion_soup[19][14] = 16'b01011_001011_00001;
        onion_soup[19][15] = 16'b01011_001011_00000;
        onion_soup[19][16] = 16'b01010_001010_00001;
        onion_soup[19][17] = 16'b01110_010000_00001;
        onion_soup[19][18] = 16'b01100_001101_00001;
        onion_soup[19][19] = 16'b01100_001100_00001;
        onion_soup[19][20] = 16'b01010_001010_00000;
        onion_soup[19][21] = 16'b01001_001001_00000;
        onion_soup[19][22] = 16'b01011_001011_00001;
        onion_soup[19][23] = 16'b01011_001011_00001;
        onion_soup[19][24] = 16'b01100_001100_00001;
        onion_soup[19][25] = 16'b10110_011101_00101;
        onion_soup[19][26] = 16'b10011_011000_00100;
        onion_soup[19][27] = 16'b11111_101011_10101;
        onion_soup[19][28] = 16'b11111_101011_10101;
        onion_soup[19][29] = 16'b11111_101011_10101;
        onion_soup[19][30] = 16'b11111_101011_10101;
        onion_soup[19][31] = 16'b11111_101011_10101;
        onion_soup[20][0] = 16'b11111_101011_10101;
        onion_soup[20][1] = 16'b11111_101011_10101;
        onion_soup[20][2] = 16'b11111_101011_10101;
        onion_soup[20][3] = 16'b11111_101011_10101;
        onion_soup[20][4] = 16'b11111_101011_10101;
        onion_soup[20][5] = 16'b11000_100010_01000;
        onion_soup[20][6] = 16'b01101_010000_00010;
        onion_soup[20][7] = 16'b10011_011010_00101;
        onion_soup[20][8] = 16'b01110_010000_00010;
        onion_soup[20][9] = 16'b01111_010010_00010;
        onion_soup[20][10] = 16'b01101_001110_00001;
        onion_soup[20][11] = 16'b10000_010010_00010;
        onion_soup[20][12] = 16'b01101_001111_00001;
        onion_soup[20][13] = 16'b01110_010000_00001;
        onion_soup[20][14] = 16'b01001_001001_00000;
        onion_soup[20][15] = 16'b01011_001100_00001;
        onion_soup[20][16] = 16'b01011_001100_00001;
        onion_soup[20][17] = 16'b01101_001110_00001;
        onion_soup[20][18] = 16'b01100_001110_00001;
        onion_soup[20][19] = 16'b01101_001111_00001;
        onion_soup[20][20] = 16'b01110_001111_00001;
        onion_soup[20][21] = 16'b01111_010001_00010;
        onion_soup[20][22] = 16'b10000_010011_00010;
        onion_soup[20][23] = 16'b01110_010000_00010;
        onion_soup[20][24] = 16'b10011_011000_00100;
        onion_soup[20][25] = 16'b10010_010110_00011;
        onion_soup[20][26] = 16'b11000_100010_00111;
        onion_soup[20][27] = 16'b11111_101011_10101;
        onion_soup[20][28] = 16'b11111_101011_10101;
        onion_soup[20][29] = 16'b11111_101011_10101;
        onion_soup[20][30] = 16'b11111_101011_10101;
        onion_soup[20][31] = 16'b11111_101011_10101;
        onion_soup[21][0] = 16'b11111_101011_10101;
        onion_soup[21][1] = 16'b11111_101011_10101;
        onion_soup[21][2] = 16'b11111_101011_10101;
        onion_soup[21][3] = 16'b11111_101011_10101;
        onion_soup[21][4] = 16'b11111_101011_10101;
        onion_soup[21][5] = 16'b11111_101011_10101;
        onion_soup[21][6] = 16'b10011_011001_00100;
        onion_soup[21][7] = 16'b10000_010100_00011;
        onion_soup[21][8] = 16'b10000_010011_00011;
        onion_soup[21][9] = 16'b10110_011101_00110;
        onion_soup[21][10] = 16'b10001_010100_00011;
        onion_soup[21][11] = 16'b10000_010011_00010;
        onion_soup[21][12] = 16'b10100_011011_00101;
        onion_soup[21][13] = 16'b10000_010100_00011;
        onion_soup[21][14] = 16'b10000_010011_00011;
        onion_soup[21][15] = 16'b10111_011110_00110;
        onion_soup[21][16] = 16'b10100_011011_00101;
        onion_soup[21][17] = 16'b10001_010110_00011;
        onion_soup[21][18] = 16'b10101_011100_00101;
        onion_soup[21][19] = 16'b10010_010110_00100;
        onion_soup[21][20] = 16'b10001_010101_00011;
        onion_soup[21][21] = 16'b10101_011011_00101;
        onion_soup[21][22] = 16'b10110_011101_00110;
        onion_soup[21][23] = 16'b10100_011001_00100;
        onion_soup[21][24] = 16'b10001_010110_00011;
        onion_soup[21][25] = 16'b10101_011101_00110;
        onion_soup[21][26] = 16'b10011_011100_00111;
        onion_soup[21][27] = 16'b11111_101011_10101;
        onion_soup[21][28] = 16'b11111_101011_10101;
        onion_soup[21][29] = 16'b11111_101011_10101;
        onion_soup[21][30] = 16'b11111_101011_10101;
        onion_soup[21][31] = 16'b11111_101011_10101;
        onion_soup[22][0] = 16'b11111_101011_10101;
        onion_soup[22][1] = 16'b11111_101011_10101;
        onion_soup[22][2] = 16'b11111_101011_10101;
        onion_soup[22][3] = 16'b11111_101011_10101;
        onion_soup[22][4] = 16'b11111_101011_10101;
        onion_soup[22][5] = 16'b11111_101011_10101;
        onion_soup[22][6] = 16'b11111_101011_10101;
        onion_soup[22][7] = 16'b11111_101011_10101;
        onion_soup[22][8] = 16'b10011_011001_00100;
        onion_soup[22][9] = 16'b01111_010010_00010;
        onion_soup[22][10] = 16'b10100_011010_00100;
        onion_soup[22][11] = 16'b10100_011001_00100;
        onion_soup[22][12] = 16'b10011_011000_00100;
        onion_soup[22][13] = 16'b10100_011001_00100;
        onion_soup[22][14] = 16'b11000_100010_01000;
        onion_soup[22][15] = 16'b10101_011011_00101;
        onion_soup[22][16] = 16'b11000_100010_01000;
        onion_soup[22][17] = 16'b11010_100111_01010;
        onion_soup[22][18] = 16'b10001_010100_00010;
        onion_soup[22][19] = 16'b11000_100011_01000;
        onion_soup[22][20] = 16'b10110_011111_00110;
        onion_soup[22][21] = 16'b10001_010101_00011;
        onion_soup[22][22] = 16'b10010_010110_00011;
        onion_soup[22][23] = 16'b10111_100000_00111;
        onion_soup[22][24] = 16'b11111_101011_10101;
        onion_soup[22][25] = 16'b11111_101011_10101;
        onion_soup[22][26] = 16'b11111_101011_10101;
        onion_soup[22][27] = 16'b11111_101011_10101;
        onion_soup[22][28] = 16'b11111_101011_10101;
        onion_soup[22][29] = 16'b11111_101011_10101;
        onion_soup[22][30] = 16'b11111_101011_10101;
        onion_soup[22][31] = 16'b11111_101011_10101;
        onion_soup[23][0] = 16'b11111_101011_10101;
        onion_soup[23][1] = 16'b11111_101011_10101;
        onion_soup[23][2] = 16'b11111_101011_10101;
        onion_soup[23][3] = 16'b11111_101011_10101;
        onion_soup[23][4] = 16'b11111_101011_10101;
        onion_soup[23][5] = 16'b11111_101011_10101;
        onion_soup[23][6] = 16'b11111_101011_10101;
        onion_soup[23][7] = 16'b11111_101011_10101;
        onion_soup[23][8] = 16'b11111_101011_10101;
        onion_soup[23][9] = 16'b11111_101011_10101;
        onion_soup[23][10] = 16'b11010_101010_01101;
        onion_soup[23][11] = 16'b11000_100100_01010;
        onion_soup[23][12] = 16'b01110_010000_00010;
        onion_soup[23][13] = 16'b10010_010110_00011;
        onion_soup[23][14] = 16'b10011_011000_00100;
        onion_soup[23][15] = 16'b10101_011100_00101;
        onion_soup[23][16] = 16'b10010_010111_00100;
        onion_soup[23][17] = 16'b10011_011000_00100;
        onion_soup[23][18] = 16'b11001_100011_00111;
        onion_soup[23][19] = 16'b10101_011011_00100;
        onion_soup[23][20] = 16'b10011_010111_00100;
        onion_soup[23][21] = 16'b11010_101011_01110;
        onion_soup[23][22] = 16'b11000_100100_01010;
        onion_soup[23][23] = 16'b11111_101011_10101;
        onion_soup[23][24] = 16'b11111_101011_10101;
        onion_soup[23][25] = 16'b11111_101011_10101;
        onion_soup[23][26] = 16'b11111_101011_10101;
        onion_soup[23][27] = 16'b11111_101011_10101;
        onion_soup[23][28] = 16'b11111_101011_10101;
        onion_soup[23][29] = 16'b11111_101011_10101;
        onion_soup[23][30] = 16'b11111_101011_10101;
        onion_soup[23][31] = 16'b11111_101011_10101;
        onion_soup[24][0] = 16'b11111_101011_10101;
        onion_soup[24][1] = 16'b11111_101011_10101;
        onion_soup[24][2] = 16'b11111_101011_10101;
        onion_soup[24][3] = 16'b11111_101011_10101;
        onion_soup[24][4] = 16'b11111_101011_10101;
        onion_soup[24][5] = 16'b11111_101011_10101;
        onion_soup[24][6] = 16'b11111_101011_10101;
        onion_soup[24][7] = 16'b11111_101011_10101;
        onion_soup[24][8] = 16'b11111_101011_10101;
        onion_soup[24][9] = 16'b11111_101011_10101;
        onion_soup[24][10] = 16'b11111_101011_10101;
        onion_soup[24][11] = 16'b11111_101011_10101;
        onion_soup[24][12] = 16'b11111_101011_10101;
        onion_soup[24][13] = 16'b11111_101011_10101;
        onion_soup[24][14] = 16'b11111_101011_10101;
        onion_soup[24][15] = 16'b11111_101011_10101;
        onion_soup[24][16] = 16'b11111_101011_10101;
        onion_soup[24][17] = 16'b11111_101011_10101;
        onion_soup[24][18] = 16'b11111_101011_10101;
        onion_soup[24][19] = 16'b11111_101011_10101;
        onion_soup[24][20] = 16'b11111_101011_10101;
        onion_soup[24][21] = 16'b11111_101011_10101;
        onion_soup[24][22] = 16'b11111_101011_10101;
        onion_soup[24][23] = 16'b11111_101011_10101;
        onion_soup[24][24] = 16'b11111_101011_10101;
        onion_soup[24][25] = 16'b11111_101011_10101;
        onion_soup[24][26] = 16'b11111_101011_10101;
        onion_soup[24][27] = 16'b11111_101011_10101;
        onion_soup[24][28] = 16'b11111_101011_10101;
        onion_soup[24][29] = 16'b11111_101011_10101;
        onion_soup[24][30] = 16'b11111_101011_10101;
        onion_soup[24][31] = 16'b11111_101011_10101;
        onion_soup[25][0] = 16'b11111_101011_10101;
        onion_soup[25][1] = 16'b11111_101011_10101;
        onion_soup[25][2] = 16'b11111_101011_10101;
        onion_soup[25][3] = 16'b11111_101011_10101;
        onion_soup[25][4] = 16'b11111_101011_10101;
        onion_soup[25][5] = 16'b11111_101011_10101;
        onion_soup[25][6] = 16'b11111_101011_10101;
        onion_soup[25][7] = 16'b11111_101011_10101;
        onion_soup[25][8] = 16'b11111_101011_10101;
        onion_soup[25][9] = 16'b11111_101011_10101;
        onion_soup[25][10] = 16'b11111_101011_10101;
        onion_soup[25][11] = 16'b11111_101011_10101;
        onion_soup[25][12] = 16'b11111_101011_10101;
        onion_soup[25][13] = 16'b11111_101011_10101;
        onion_soup[25][14] = 16'b11111_101011_10101;
        onion_soup[25][15] = 16'b11111_101011_10101;
        onion_soup[25][16] = 16'b11111_101011_10101;
        onion_soup[25][17] = 16'b11111_101011_10101;
        onion_soup[25][18] = 16'b11111_101011_10101;
        onion_soup[25][19] = 16'b11111_101011_10101;
        onion_soup[25][20] = 16'b11111_101011_10101;
        onion_soup[25][21] = 16'b11111_101011_10101;
        onion_soup[25][22] = 16'b11111_101011_10101;
        onion_soup[25][23] = 16'b11111_101011_10101;
        onion_soup[25][24] = 16'b11111_101011_10101;
        onion_soup[25][25] = 16'b11111_101011_10101;
        onion_soup[25][26] = 16'b11111_101011_10101;
        onion_soup[25][27] = 16'b11111_101011_10101;
        onion_soup[25][28] = 16'b11111_101011_10101;
        onion_soup[25][29] = 16'b11111_101011_10101;
        onion_soup[25][30] = 16'b11111_101011_10101;
        onion_soup[25][31] = 16'b11111_101011_10101;
        onion_soup[26][0] = 16'b11111_101011_10101;
        onion_soup[26][1] = 16'b11111_101011_10101;
        onion_soup[26][2] = 16'b11111_101011_10101;
        onion_soup[26][3] = 16'b11111_101011_10101;
        onion_soup[26][4] = 16'b11111_101011_10101;
        onion_soup[26][5] = 16'b11111_101011_10101;
        onion_soup[26][6] = 16'b11111_101011_10101;
        onion_soup[26][7] = 16'b11111_101011_10101;
        onion_soup[26][8] = 16'b11111_101011_10101;
        onion_soup[26][9] = 16'b11111_101011_10101;
        onion_soup[26][10] = 16'b11111_101011_10101;
        onion_soup[26][11] = 16'b11111_101011_10101;
        onion_soup[26][12] = 16'b11111_101011_10101;
        onion_soup[26][13] = 16'b11111_101011_10101;
        onion_soup[26][14] = 16'b11111_101011_10101;
        onion_soup[26][15] = 16'b11111_101011_10101;
        onion_soup[26][16] = 16'b11111_101011_10101;
        onion_soup[26][17] = 16'b11111_101011_10101;
        onion_soup[26][18] = 16'b11111_101011_10101;
        onion_soup[26][19] = 16'b11111_101011_10101;
        onion_soup[26][20] = 16'b11111_101011_10101;
        onion_soup[26][21] = 16'b11111_101011_10101;
        onion_soup[26][22] = 16'b11111_101011_10101;
        onion_soup[26][23] = 16'b11111_101011_10101;
        onion_soup[26][24] = 16'b11111_101011_10101;
        onion_soup[26][25] = 16'b11111_101011_10101;
        onion_soup[26][26] = 16'b11111_101011_10101;
        onion_soup[26][27] = 16'b11111_101011_10101;
        onion_soup[26][28] = 16'b11111_101011_10101;
        onion_soup[26][29] = 16'b11111_101011_10101;
        onion_soup[26][30] = 16'b11111_101011_10101;
        onion_soup[26][31] = 16'b11111_101011_10101;
        onion_soup[27][0] = 16'b11111_101011_10101;
        onion_soup[27][1] = 16'b11111_101011_10101;
        onion_soup[27][2] = 16'b11111_101011_10101;
        onion_soup[27][3] = 16'b11111_101011_10101;
        onion_soup[27][4] = 16'b11111_101011_10101;
        onion_soup[27][5] = 16'b11111_101011_10101;
        onion_soup[27][6] = 16'b11111_101011_10101;
        onion_soup[27][7] = 16'b11111_101011_10101;
        onion_soup[27][8] = 16'b11111_101011_10101;
        onion_soup[27][9] = 16'b11111_101011_10101;
        onion_soup[27][10] = 16'b11111_101011_10101;
        onion_soup[27][11] = 16'b11111_101011_10101;
        onion_soup[27][12] = 16'b11111_101011_10101;
        onion_soup[27][13] = 16'b11111_101011_10101;
        onion_soup[27][14] = 16'b11111_101011_10101;
        onion_soup[27][15] = 16'b11111_101011_10101;
        onion_soup[27][16] = 16'b11111_101011_10101;
        onion_soup[27][17] = 16'b11111_101011_10101;
        onion_soup[27][18] = 16'b11111_101011_10101;
        onion_soup[27][19] = 16'b11111_101011_10101;
        onion_soup[27][20] = 16'b11111_101011_10101;
        onion_soup[27][21] = 16'b11111_101011_10101;
        onion_soup[27][22] = 16'b11111_101011_10101;
        onion_soup[27][23] = 16'b11111_101011_10101;
        onion_soup[27][24] = 16'b11111_101011_10101;
        onion_soup[27][25] = 16'b11111_101011_10101;
        onion_soup[27][26] = 16'b11111_101011_10101;
        onion_soup[27][27] = 16'b11111_101011_10101;
        onion_soup[27][28] = 16'b11111_101011_10101;
        onion_soup[27][29] = 16'b11111_101011_10101;
        onion_soup[27][30] = 16'b11111_101011_10101;
        onion_soup[27][31] = 16'b11111_101011_10101;
        onion_soup[28][0] = 16'b11111_101011_10101;
        onion_soup[28][1] = 16'b11111_101011_10101;
        onion_soup[28][2] = 16'b11111_101011_10101;
        onion_soup[28][3] = 16'b11111_101011_10101;
        onion_soup[28][4] = 16'b11111_101011_10101;
        onion_soup[28][5] = 16'b11111_101011_10101;
        onion_soup[28][6] = 16'b11111_101011_10101;
        onion_soup[28][7] = 16'b11111_101011_10101;
        onion_soup[28][8] = 16'b11111_101011_10101;
        onion_soup[28][9] = 16'b11111_101011_10101;
        onion_soup[28][10] = 16'b11111_101011_10101;
        onion_soup[28][11] = 16'b11111_101011_10101;
        onion_soup[28][12] = 16'b11111_101011_10101;
        onion_soup[28][13] = 16'b11111_101011_10101;
        onion_soup[28][14] = 16'b11111_101011_10101;
        onion_soup[28][15] = 16'b11111_101011_10101;
        onion_soup[28][16] = 16'b11111_101011_10101;
        onion_soup[28][17] = 16'b11111_101011_10101;
        onion_soup[28][18] = 16'b11111_101011_10101;
        onion_soup[28][19] = 16'b11111_101011_10101;
        onion_soup[28][20] = 16'b11111_101011_10101;
        onion_soup[28][21] = 16'b11111_101011_10101;
        onion_soup[28][22] = 16'b11111_101011_10101;
        onion_soup[28][23] = 16'b11111_101011_10101;
        onion_soup[28][24] = 16'b11111_101011_10101;
        onion_soup[28][25] = 16'b11111_101011_10101;
        onion_soup[28][26] = 16'b11111_101011_10101;
        onion_soup[28][27] = 16'b11111_101011_10101;
        onion_soup[28][28] = 16'b11111_101011_10101;
        onion_soup[28][29] = 16'b11111_101011_10101;
        onion_soup[28][30] = 16'b11111_101011_10101;
        onion_soup[28][31] = 16'b11111_101011_10101;
        onion_soup[29][0] = 16'b11111_101011_10101;
        onion_soup[29][1] = 16'b11111_101011_10101;
        onion_soup[29][2] = 16'b11111_101011_10101;
        onion_soup[29][3] = 16'b11111_101011_10101;
        onion_soup[29][4] = 16'b11111_101011_10101;
        onion_soup[29][5] = 16'b11111_101011_10101;
        onion_soup[29][6] = 16'b11111_101011_10101;
        onion_soup[29][7] = 16'b11111_101011_10101;
        onion_soup[29][8] = 16'b11111_101011_10101;
        onion_soup[29][9] = 16'b11111_101011_10101;
        onion_soup[29][10] = 16'b11111_101011_10101;
        onion_soup[29][11] = 16'b11111_101011_10101;
        onion_soup[29][12] = 16'b11111_101011_10101;
        onion_soup[29][13] = 16'b11111_101011_10101;
        onion_soup[29][14] = 16'b11111_101011_10101;
        onion_soup[29][15] = 16'b11111_101011_10101;
        onion_soup[29][16] = 16'b11111_101011_10101;
        onion_soup[29][17] = 16'b11111_101011_10101;
        onion_soup[29][18] = 16'b11111_101011_10101;
        onion_soup[29][19] = 16'b11111_101011_10101;
        onion_soup[29][20] = 16'b11111_101011_10101;
        onion_soup[29][21] = 16'b11111_101011_10101;
        onion_soup[29][22] = 16'b11111_101011_10101;
        onion_soup[29][23] = 16'b11111_101011_10101;
        onion_soup[29][24] = 16'b11111_101011_10101;
        onion_soup[29][25] = 16'b11111_101011_10101;
        onion_soup[29][26] = 16'b11111_101011_10101;
        onion_soup[29][27] = 16'b11111_101011_10101;
        onion_soup[29][28] = 16'b11111_101011_10101;
        onion_soup[29][29] = 16'b11111_101011_10101;
        onion_soup[29][30] = 16'b11111_101011_10101;
        onion_soup[29][31] = 16'b11111_101011_10101;
        onion_soup[30][0] = 16'b11111_101011_10101;
        onion_soup[30][1] = 16'b11111_101011_10101;
        onion_soup[30][2] = 16'b11111_101011_10101;
        onion_soup[30][3] = 16'b11111_101011_10101;
        onion_soup[30][4] = 16'b11111_101011_10101;
        onion_soup[30][5] = 16'b11111_101011_10101;
        onion_soup[30][6] = 16'b11111_101011_10101;
        onion_soup[30][7] = 16'b11111_101011_10101;
        onion_soup[30][8] = 16'b11111_101011_10101;
        onion_soup[30][9] = 16'b11111_101011_10101;
        onion_soup[30][10] = 16'b11111_101011_10101;
        onion_soup[30][11] = 16'b11111_101011_10101;
        onion_soup[30][12] = 16'b11111_101011_10101;
        onion_soup[30][13] = 16'b11111_101011_10101;
        onion_soup[30][14] = 16'b11111_101011_10101;
        onion_soup[30][15] = 16'b11111_101011_10101;
        onion_soup[30][16] = 16'b11111_101011_10101;
        onion_soup[30][17] = 16'b11111_101011_10101;
        onion_soup[30][18] = 16'b11111_101011_10101;
        onion_soup[30][19] = 16'b11111_101011_10101;
        onion_soup[30][20] = 16'b11111_101011_10101;
        onion_soup[30][21] = 16'b11111_101011_10101;
        onion_soup[30][22] = 16'b11111_101011_10101;
        onion_soup[30][23] = 16'b11111_101011_10101;
        onion_soup[30][24] = 16'b11111_101011_10101;
        onion_soup[30][25] = 16'b11111_101011_10101;
        onion_soup[30][26] = 16'b11111_101011_10101;
        onion_soup[30][27] = 16'b11111_101011_10101;
        onion_soup[30][28] = 16'b11111_101011_10101;
        onion_soup[30][29] = 16'b11111_101011_10101;
        onion_soup[30][30] = 16'b11111_101011_10101;
        onion_soup[30][31] = 16'b11111_101011_10101;
        onion_soup[31][0] = 16'b11111_101011_10101;
        onion_soup[31][1] = 16'b11111_101011_10101;
        onion_soup[31][2] = 16'b11111_101011_10101;
        onion_soup[31][3] = 16'b11111_101011_10101;
        onion_soup[31][4] = 16'b11111_101011_10101;
        onion_soup[31][5] = 16'b11111_101011_10101;
        onion_soup[31][6] = 16'b11111_101011_10101;
        onion_soup[31][7] = 16'b11111_101011_10101;
        onion_soup[31][8] = 16'b11111_101011_10101;
        onion_soup[31][9] = 16'b11111_101011_10101;
        onion_soup[31][10] = 16'b11111_101011_10101;
        onion_soup[31][11] = 16'b11111_101011_10101;
        onion_soup[31][12] = 16'b11111_101011_10101;
        onion_soup[31][13] = 16'b11111_101011_10101;
        onion_soup[31][14] = 16'b11111_101011_10101;
        onion_soup[31][15] = 16'b11111_101011_10101;
        onion_soup[31][16] = 16'b11111_101011_10101;
        onion_soup[31][17] = 16'b11111_101011_10101;
        onion_soup[31][18] = 16'b11111_101011_10101;
        onion_soup[31][19] = 16'b11111_101011_10101;
        onion_soup[31][20] = 16'b11111_101011_10101;
        onion_soup[31][21] = 16'b11111_101011_10101;
        onion_soup[31][22] = 16'b11111_101011_10101;
        onion_soup[31][23] = 16'b11111_101011_10101;
        onion_soup[31][24] = 16'b11111_101011_10101;
        onion_soup[31][25] = 16'b11111_101011_10101;
        onion_soup[31][26] = 16'b11111_101011_10101;
        onion_soup[31][27] = 16'b11111_101011_10101;
        onion_soup[31][28] = 16'b11111_101011_10101;
        onion_soup[31][29] = 16'b11111_101011_10101;
        onion_soup[31][30] = 16'b11111_101011_10101;
        onion_soup[31][31] = 16'b11111_101011_10101;



        
        tomato_soup[0][0] = 16'b10111_111111_10101;
        tomato_soup[0][1] = 16'b10111_111111_10101;
        tomato_soup[0][2] = 16'b10111_111111_10101;
        tomato_soup[0][3] = 16'b10111_111111_10101;
        tomato_soup[0][4] = 16'b10111_111111_10101;
        tomato_soup[0][5] = 16'b10111_111111_10101;
        tomato_soup[0][6] = 16'b10111_111111_10101;
        tomato_soup[0][7] = 16'b10111_111111_10101;
        tomato_soup[0][8] = 16'b10111_111111_10101;
        tomato_soup[0][9] = 16'b10111_111111_10101;
        tomato_soup[0][10] = 16'b10111_111111_10101;
        tomato_soup[0][11] = 16'b10111_111111_10101;
        tomato_soup[0][12] = 16'b10111_111111_10101;
        tomato_soup[0][13] = 16'b10111_111111_10101;
        tomato_soup[0][14] = 16'b10111_111111_10101;
        tomato_soup[0][15] = 16'b10111_111111_10101;
        tomato_soup[0][16] = 16'b10111_111111_10101;
        tomato_soup[0][17] = 16'b10111_111111_10101;
        tomato_soup[0][18] = 16'b10111_111111_10101;
        tomato_soup[0][19] = 16'b10111_111111_10101;
        tomato_soup[0][20] = 16'b10111_111111_10101;
        tomato_soup[0][21] = 16'b10111_111111_10101;
        tomato_soup[0][22] = 16'b10111_111111_10101;
        tomato_soup[0][23] = 16'b10111_111111_10101;
        tomato_soup[0][24] = 16'b10111_111111_10101;
        tomato_soup[0][25] = 16'b10111_111111_10101;
        tomato_soup[0][26] = 16'b10111_111111_10101;
        tomato_soup[0][27] = 16'b10111_111111_10101;
        tomato_soup[0][28] = 16'b10111_111111_10101;
        tomato_soup[0][29] = 16'b10111_111111_10101;
        tomato_soup[0][30] = 16'b10111_111111_10101;
        tomato_soup[0][31] = 16'b10111_111111_10101;
        tomato_soup[1][0] = 16'b10111_111111_10101;
        tomato_soup[1][1] = 16'b10111_111111_10101;
        tomato_soup[1][2] = 16'b10111_111111_10101;
        tomato_soup[1][3] = 16'b10111_111111_10101;
        tomato_soup[1][4] = 16'b10111_111111_10101;
        tomato_soup[1][5] = 16'b10111_111111_10101;
        tomato_soup[1][6] = 16'b10111_111111_10101;
        tomato_soup[1][7] = 16'b10111_111111_10101;
        tomato_soup[1][8] = 16'b10111_111111_10101;
        tomato_soup[1][9] = 16'b10111_111111_10101;
        tomato_soup[1][10] = 16'b10111_111111_10101;
        tomato_soup[1][11] = 16'b10111_111111_10101;
        tomato_soup[1][12] = 16'b10111_111111_10101;
        tomato_soup[1][13] = 16'b10111_111111_10101;
        tomato_soup[1][14] = 16'b10111_111111_10101;
        tomato_soup[1][15] = 16'b10111_111111_10101;
        tomato_soup[1][16] = 16'b10111_111111_10101;
        tomato_soup[1][17] = 16'b10111_111111_10101;
        tomato_soup[1][18] = 16'b10111_111111_10101;
        tomato_soup[1][19] = 16'b10111_111111_10101;
        tomato_soup[1][20] = 16'b10111_111111_10101;
        tomato_soup[1][21] = 16'b10111_111111_10101;
        tomato_soup[1][22] = 16'b10111_111111_10101;
        tomato_soup[1][23] = 16'b10111_111111_10101;
        tomato_soup[1][24] = 16'b10111_111111_10101;
        tomato_soup[1][25] = 16'b10111_111111_10101;
        tomato_soup[1][26] = 16'b10111_111111_10101;
        tomato_soup[1][27] = 16'b10111_111111_10101;
        tomato_soup[1][28] = 16'b10111_111111_10101;
        tomato_soup[1][29] = 16'b10111_111111_10101;
        tomato_soup[1][30] = 16'b10111_111111_10101;
        tomato_soup[1][31] = 16'b10111_111111_10101;
        tomato_soup[2][0] = 16'b10111_111111_10101;
        tomato_soup[2][1] = 16'b10111_111111_10101;
        tomato_soup[2][2] = 16'b10111_111111_10101;
        tomato_soup[2][3] = 16'b10111_111111_10101;
        tomato_soup[2][4] = 16'b10111_111111_10101;
        tomato_soup[2][5] = 16'b10111_111111_10101;
        tomato_soup[2][6] = 16'b10111_111111_10101;
        tomato_soup[2][7] = 16'b10111_111111_10101;
        tomato_soup[2][8] = 16'b10111_111111_10101;
        tomato_soup[2][9] = 16'b10111_111111_10101;
        tomato_soup[2][10] = 16'b10111_111111_10101;
        tomato_soup[2][11] = 16'b10111_111111_10101;
        tomato_soup[2][12] = 16'b10111_111111_10101;
        tomato_soup[2][13] = 16'b10111_111111_10101;
        tomato_soup[2][14] = 16'b10111_111111_10101;
        tomato_soup[2][15] = 16'b10111_111111_10101;
        tomato_soup[2][16] = 16'b10111_111111_10101;
        tomato_soup[2][17] = 16'b10111_111111_10101;
        tomato_soup[2][18] = 16'b10111_111111_10101;
        tomato_soup[2][19] = 16'b10111_111111_10101;
        tomato_soup[2][20] = 16'b10111_111111_10101;
        tomato_soup[2][21] = 16'b10111_111111_10101;
        tomato_soup[2][22] = 16'b10111_111111_10101;
        tomato_soup[2][23] = 16'b10111_111111_10101;
        tomato_soup[2][24] = 16'b10111_111111_10101;
        tomato_soup[2][25] = 16'b10111_111111_10101;
        tomato_soup[2][26] = 16'b10111_111111_10101;
        tomato_soup[2][27] = 16'b10111_111111_10101;
        tomato_soup[2][28] = 16'b10111_111111_10101;
        tomato_soup[2][29] = 16'b10111_111111_10101;
        tomato_soup[2][30] = 16'b10111_111111_10101;
        tomato_soup[2][31] = 16'b10111_111111_10101;
        tomato_soup[3][0] = 16'b10111_111111_10101;
        tomato_soup[3][1] = 16'b10111_111111_10101;
        tomato_soup[3][2] = 16'b10111_111111_10101;
        tomato_soup[3][3] = 16'b10111_111111_10101;
        tomato_soup[3][4] = 16'b10111_111111_10101;
        tomato_soup[3][5] = 16'b10111_111111_10101;
        tomato_soup[3][6] = 16'b10111_111111_10101;
        tomato_soup[3][7] = 16'b10111_111111_10101;
        tomato_soup[3][8] = 16'b10111_111111_10101;
        tomato_soup[3][9] = 16'b10111_111111_10101;
        tomato_soup[3][10] = 16'b10111_111111_10101;
        tomato_soup[3][11] = 16'b10111_111111_10101;
        tomato_soup[3][12] = 16'b10111_111111_10101;
        tomato_soup[3][13] = 16'b10111_111111_10101;
        tomato_soup[3][14] = 16'b10111_111111_10101;
        tomato_soup[3][15] = 16'b10111_111111_10101;
        tomato_soup[3][16] = 16'b10111_111111_10101;
        tomato_soup[3][17] = 16'b10111_111111_10101;
        tomato_soup[3][18] = 16'b10111_111111_10101;
        tomato_soup[3][19] = 16'b10111_111111_10101;
        tomato_soup[3][20] = 16'b10111_111111_10101;
        tomato_soup[3][21] = 16'b10111_111111_10101;
        tomato_soup[3][22] = 16'b10111_111111_10101;
        tomato_soup[3][23] = 16'b10111_111111_10101;
        tomato_soup[3][24] = 16'b10111_111111_10101;
        tomato_soup[3][25] = 16'b10111_111111_10101;
        tomato_soup[3][26] = 16'b10111_111111_10101;
        tomato_soup[3][27] = 16'b10111_111111_10101;
        tomato_soup[3][28] = 16'b10111_111111_10101;
        tomato_soup[3][29] = 16'b10111_111111_10101;
        tomato_soup[3][30] = 16'b10111_111111_10101;
        tomato_soup[3][31] = 16'b10111_111111_10101;
        tomato_soup[4][0] = 16'b10111_111111_10101;
        tomato_soup[4][1] = 16'b10111_111111_10101;
        tomato_soup[4][2] = 16'b10111_111111_10101;
        tomato_soup[4][3] = 16'b10111_111111_10101;
        tomato_soup[4][4] = 16'b10111_111111_10101;
        tomato_soup[4][5] = 16'b10111_111111_10101;
        tomato_soup[4][6] = 16'b10111_111111_10101;
        tomato_soup[4][7] = 16'b10111_111111_10101;
        tomato_soup[4][8] = 16'b10111_111111_10101;
        tomato_soup[4][9] = 16'b10111_111111_10101;
        tomato_soup[4][10] = 16'b10111_111111_10101;
        tomato_soup[4][11] = 16'b11001_101000_01100;
        tomato_soup[4][12] = 16'b11001_101000_01100;
        tomato_soup[4][13] = 16'b11000_100111_01100;
        tomato_soup[4][14] = 16'b11000_101000_01100;
        tomato_soup[4][15] = 16'b11000_101000_01100;
        tomato_soup[4][16] = 16'b11000_101000_01100;
        tomato_soup[4][17] = 16'b11001_101000_01100;
        tomato_soup[4][18] = 16'b11000_101000_01100;
        tomato_soup[4][19] = 16'b11001_101001_01101;
        tomato_soup[4][20] = 16'b10111_111111_10101;
        tomato_soup[4][21] = 16'b10111_111111_10101;
        tomato_soup[4][22] = 16'b10111_111111_10101;
        tomato_soup[4][23] = 16'b10111_111111_10101;
        tomato_soup[4][24] = 16'b10111_111111_10101;
        tomato_soup[4][25] = 16'b10111_111111_10101;
        tomato_soup[4][26] = 16'b10111_111111_10101;
        tomato_soup[4][27] = 16'b10111_111111_10101;
        tomato_soup[4][28] = 16'b10111_111111_10101;
        tomato_soup[4][29] = 16'b10111_111111_10101;
        tomato_soup[4][30] = 16'b10111_111111_10101;
        tomato_soup[4][31] = 16'b10111_111111_10101;
        tomato_soup[5][0] = 16'b10111_111111_10101;
        tomato_soup[5][1] = 16'b10111_111111_10101;
        tomato_soup[5][2] = 16'b10111_111111_10101;
        tomato_soup[5][3] = 16'b10111_111111_10101;
        tomato_soup[5][4] = 16'b10111_111111_10101;
        tomato_soup[5][5] = 16'b10111_111111_10101;
        tomato_soup[5][6] = 16'b10111_111111_10101;
        tomato_soup[5][7] = 16'b10111_111111_10101;
        tomato_soup[5][8] = 16'b10111_111111_10101;
        tomato_soup[5][9] = 16'b11001_101001_01101;
        tomato_soup[5][10] = 16'b11001_101000_01101;
        tomato_soup[5][11] = 16'b11001_101001_01101;
        tomato_soup[5][12] = 16'b11001_101010_01110;
        tomato_soup[5][13] = 16'b11001_101010_01101;
        tomato_soup[5][14] = 16'b11001_101010_01110;
        tomato_soup[5][15] = 16'b11010_101100_01111;
        tomato_soup[5][16] = 16'b11001_101010_01110;
        tomato_soup[5][17] = 16'b11010_101011_01110;
        tomato_soup[5][18] = 16'b11010_101011_01110;
        tomato_soup[5][19] = 16'b11001_101011_01110;
        tomato_soup[5][20] = 16'b11001_101001_01101;
        tomato_soup[5][21] = 16'b11001_101001_01101;
        tomato_soup[5][22] = 16'b10111_111111_10101;
        tomato_soup[5][23] = 16'b10111_111111_10101;
        tomato_soup[5][24] = 16'b10111_111111_10101;
        tomato_soup[5][25] = 16'b10111_111111_10101;
        tomato_soup[5][26] = 16'b10111_111111_10101;
        tomato_soup[5][27] = 16'b10111_111111_10101;
        tomato_soup[5][28] = 16'b10111_111111_10101;
        tomato_soup[5][29] = 16'b10111_111111_10101;
        tomato_soup[5][30] = 16'b10111_111111_10101;
        tomato_soup[5][31] = 16'b10111_111111_10101;
        tomato_soup[6][0] = 16'b10111_111111_10101;
        tomato_soup[6][1] = 16'b10111_111111_10101;
        tomato_soup[6][2] = 16'b10111_111111_10101;
        tomato_soup[6][3] = 16'b10111_111111_10101;
        tomato_soup[6][4] = 16'b10111_111111_10101;
        tomato_soup[6][5] = 16'b10111_111111_10101;
        tomato_soup[6][6] = 16'b10111_111111_10101;
        tomato_soup[6][7] = 16'b11001_101001_01101;
        tomato_soup[6][8] = 16'b11001_101001_01101;
        tomato_soup[6][9] = 16'b11001_101010_01110;
        tomato_soup[6][10] = 16'b11010_101011_01110;
        tomato_soup[6][11] = 16'b11010_101011_01110;
        tomato_soup[6][12] = 16'b11010_101011_01110;
        tomato_soup[6][13] = 16'b11001_101010_01110;
        tomato_soup[6][14] = 16'b11001_101011_01110;
        tomato_soup[6][15] = 16'b11001_101010_01101;
        tomato_soup[6][16] = 16'b11001_101010_01101;
        tomato_soup[6][17] = 16'b11001_101001_01101;
        tomato_soup[6][18] = 16'b11001_101010_01110;
        tomato_soup[6][19] = 16'b11001_101010_01110;
        tomato_soup[6][20] = 16'b11010_101011_01110;
        tomato_soup[6][21] = 16'b11001_101010_01101;
        tomato_soup[6][22] = 16'b11001_101001_01101;
        tomato_soup[6][23] = 16'b11001_101001_01101;
        tomato_soup[6][24] = 16'b10111_111111_10101;
        tomato_soup[6][25] = 16'b10111_111111_10101;
        tomato_soup[6][26] = 16'b10111_111111_10101;
        tomato_soup[6][27] = 16'b10111_111111_10101;
        tomato_soup[6][28] = 16'b10111_111111_10101;
        tomato_soup[6][29] = 16'b10111_111111_10101;
        tomato_soup[6][30] = 16'b10111_111111_10101;
        tomato_soup[6][31] = 16'b10111_111111_10101;
        tomato_soup[7][0] = 16'b10111_111111_10101;
        tomato_soup[7][1] = 16'b10111_111111_10101;
        tomato_soup[7][2] = 16'b10111_111111_10101;
        tomato_soup[7][3] = 16'b10111_111111_10101;
        tomato_soup[7][4] = 16'b10111_111111_10101;
        tomato_soup[7][5] = 16'b10111_111111_10101;
        tomato_soup[7][6] = 16'b11001_101001_01101;
        tomato_soup[7][7] = 16'b11001_101001_01101;
        tomato_soup[7][8] = 16'b11001_101010_01110;
        tomato_soup[7][9] = 16'b11001_101010_01110;
        tomato_soup[7][10] = 16'b11001_101010_01110;
        tomato_soup[7][11] = 16'b11001_101011_01110;
        tomato_soup[7][12] = 16'b11001_101010_01101;
        tomato_soup[7][13] = 16'b11001_101010_01110;
        tomato_soup[7][14] = 16'b11001_101010_01110;
        tomato_soup[7][15] = 16'b11001_101010_01101;
        tomato_soup[7][16] = 16'b11001_101010_01110;
        tomato_soup[7][17] = 16'b11010_101011_01110;
        tomato_soup[7][18] = 16'b11001_101001_01101;
        tomato_soup[7][19] = 16'b11001_101010_01101;
        tomato_soup[7][20] = 16'b11010_101100_01111;
        tomato_soup[7][21] = 16'b11010_101011_01110;
        tomato_soup[7][22] = 16'b11001_101010_01110;
        tomato_soup[7][23] = 16'b11010_101011_01110;
        tomato_soup[7][24] = 16'b11001_101010_01101;
        tomato_soup[7][25] = 16'b10111_111111_10101;
        tomato_soup[7][26] = 16'b10111_111111_10101;
        tomato_soup[7][27] = 16'b10111_111111_10101;
        tomato_soup[7][28] = 16'b10111_111111_10101;
        tomato_soup[7][29] = 16'b10111_111111_10101;
        tomato_soup[7][30] = 16'b10111_111111_10101;
        tomato_soup[7][31] = 16'b10111_111111_10101;
        tomato_soup[8][0] = 16'b10111_111111_10101;
        tomato_soup[8][1] = 16'b10111_111111_10101;
        tomato_soup[8][2] = 16'b10111_111111_10101;
        tomato_soup[8][3] = 16'b10111_111111_10101;
        tomato_soup[8][4] = 16'b10111_111111_10101;
        tomato_soup[8][5] = 16'b11001_101001_01101;
        tomato_soup[8][6] = 16'b11001_101001_01101;
        tomato_soup[8][7] = 16'b11001_101010_01110;
        tomato_soup[8][8] = 16'b11001_101010_01110;
        tomato_soup[8][9] = 16'b11001_101001_01101;
        tomato_soup[8][10] = 16'b11001_101010_01110;
        tomato_soup[8][11] = 16'b11001_101010_01101;
        tomato_soup[8][12] = 16'b11001_101001_01101;
        tomato_soup[8][13] = 16'b11001_101001_01101;
        tomato_soup[8][14] = 16'b11001_101001_01101;
        tomato_soup[8][15] = 16'b11001_101010_01110;
        tomato_soup[8][16] = 16'b11001_101001_01101;
        tomato_soup[8][17] = 16'b11001_101001_01101;
        tomato_soup[8][18] = 16'b11001_101001_01101;
        tomato_soup[8][19] = 16'b11001_101001_01101;
        tomato_soup[8][20] = 16'b11001_101010_01110;
        tomato_soup[8][21] = 16'b11001_101001_01101;
        tomato_soup[8][22] = 16'b11001_101010_01110;
        tomato_soup[8][23] = 16'b11001_101011_01110;
        tomato_soup[8][24] = 16'b11001_101010_01110;
        tomato_soup[8][25] = 16'b11001_101010_01101;
        tomato_soup[8][26] = 16'b10111_111111_10101;
        tomato_soup[8][27] = 16'b10111_111111_10101;
        tomato_soup[8][28] = 16'b10111_111111_10101;
        tomato_soup[8][29] = 16'b10111_111111_10101;
        tomato_soup[8][30] = 16'b10111_111111_10101;
        tomato_soup[8][31] = 16'b10111_111111_10101;
        tomato_soup[9][0] = 16'b10111_111111_10101;
        tomato_soup[9][1] = 16'b10111_111111_10101;
        tomato_soup[9][2] = 16'b10111_111111_10101;
        tomato_soup[9][3] = 16'b10111_111111_10101;
        tomato_soup[9][4] = 16'b10111_111111_10101;
        tomato_soup[9][5] = 16'b11001_101010_01101;
        tomato_soup[9][6] = 16'b11001_101010_01110;
        tomato_soup[9][7] = 16'b11001_101001_01101;
        tomato_soup[9][8] = 16'b11001_101001_01101;
        tomato_soup[9][9] = 16'b11001_101010_01110;
        tomato_soup[9][10] = 16'b11001_101010_01110;
        tomato_soup[9][11] = 16'b11001_101011_01110;
        tomato_soup[9][12] = 16'b11010_101101_10000;
        tomato_soup[9][13] = 16'b11011_101110_10001;
        tomato_soup[9][14] = 16'b11010_101101_10000;
        tomato_soup[9][15] = 16'b11010_101100_01111;
        tomato_soup[9][16] = 16'b11010_101101_10000;
        tomato_soup[9][17] = 16'b11011_101110_10000;
        tomato_soup[9][18] = 16'b11011_101110_10000;
        tomato_soup[9][19] = 16'b11010_101101_10000;
        tomato_soup[9][20] = 16'b11001_101010_01101;
        tomato_soup[9][21] = 16'b11001_101001_01101;
        tomato_soup[9][22] = 16'b11001_101010_01101;
        tomato_soup[9][23] = 16'b11001_101010_01101;
        tomato_soup[9][24] = 16'b11001_101010_01110;
        tomato_soup[9][25] = 16'b11001_101001_01101;
        tomato_soup[9][26] = 16'b11001_101001_01101;
        tomato_soup[9][27] = 16'b10111_111111_10101;
        tomato_soup[9][28] = 16'b10111_111111_10101;
        tomato_soup[9][29] = 16'b10111_111111_10101;
        tomato_soup[9][30] = 16'b10111_111111_10101;
        tomato_soup[9][31] = 16'b10111_111111_10101;
        tomato_soup[10][0] = 16'b10111_111111_10101;
        tomato_soup[10][1] = 16'b10111_111111_10101;
        tomato_soup[10][2] = 16'b10111_111111_10101;
        tomato_soup[10][3] = 16'b10111_111111_10101;
        tomato_soup[10][4] = 16'b11001_101001_01101;
        tomato_soup[10][5] = 16'b11001_101001_01101;
        tomato_soup[10][6] = 16'b11001_101001_01101;
        tomato_soup[10][7] = 16'b11001_101001_01101;
        tomato_soup[10][8] = 16'b11010_101101_10000;
        tomato_soup[10][9] = 16'b11011_101111_10001;
        tomato_soup[10][10] = 16'b11011_101110_10000;
        tomato_soup[10][11] = 16'b11010_101100_01111;
        tomato_soup[10][12] = 16'b11001_101001_01101;
        tomato_soup[10][13] = 16'b11000_011110_00111;
        tomato_soup[10][14] = 16'b11000_011000_00101;
        tomato_soup[10][15] = 16'b11000_011000_00101;
        tomato_soup[10][16] = 16'b11000_011010_00110;
        tomato_soup[10][17] = 16'b11000_011101_00111;
        tomato_soup[10][18] = 16'b11001_100011_01010;
        tomato_soup[10][19] = 16'b11010_101100_01111;
        tomato_soup[10][20] = 16'b11010_101100_01111;
        tomato_soup[10][21] = 16'b11010_101100_01111;
        tomato_soup[10][22] = 16'b11010_101101_10000;
        tomato_soup[10][23] = 16'b11001_101010_01101;
        tomato_soup[10][24] = 16'b11001_101001_01101;
        tomato_soup[10][25] = 16'b11001_101010_01101;
        tomato_soup[10][26] = 16'b11001_101010_01101;
        tomato_soup[10][27] = 16'b10111_111111_10101;
        tomato_soup[10][28] = 16'b10111_111111_10101;
        tomato_soup[10][29] = 16'b10111_111111_10101;
        tomato_soup[10][30] = 16'b10111_111111_10101;
        tomato_soup[10][31] = 16'b10111_111111_10101;
        tomato_soup[11][0] = 16'b10111_111111_10101;
        tomato_soup[11][1] = 16'b10111_111111_10101;
        tomato_soup[11][2] = 16'b10111_111111_10101;
        tomato_soup[11][3] = 16'b10111_111111_10101;
        tomato_soup[11][4] = 16'b11001_101001_01101;
        tomato_soup[11][5] = 16'b11001_101001_01101;
        tomato_soup[11][6] = 16'b11010_101101_10000;
        tomato_soup[11][7] = 16'b11011_101101_10000;
        tomato_soup[11][8] = 16'b11010_101101_10000;
        tomato_soup[11][9] = 16'b11000_011101_00111;
        tomato_soup[11][10] = 16'b10111_010010_00010;
        tomato_soup[11][11] = 16'b10111_001101_00001;
        tomato_soup[11][12] = 16'b10111_001100_00001;
        tomato_soup[11][13] = 16'b10111_001011_00001;
        tomato_soup[11][14] = 16'b11000_001101_00001;
        tomato_soup[11][15] = 16'b10111_001100_00001;
        tomato_soup[11][16] = 16'b10111_001100_00001;
        tomato_soup[11][17] = 16'b10111_001011_00001;
        tomato_soup[11][18] = 16'b10111_001100_00001;
        tomato_soup[11][19] = 16'b10111_001011_00001;
        tomato_soup[11][20] = 16'b10111_001011_00001;
        tomato_soup[11][21] = 16'b11000_011001_00101;
        tomato_soup[11][22] = 16'b11011_101110_10000;
        tomato_soup[11][23] = 16'b11011_110000_10010;
        tomato_soup[11][24] = 16'b11011_101111_10001;
        tomato_soup[11][25] = 16'b11001_101001_01101;
        tomato_soup[11][26] = 16'b11001_101001_01101;
        tomato_soup[11][27] = 16'b11001_101000_01100;
        tomato_soup[11][28] = 16'b10111_111111_10101;
        tomato_soup[11][29] = 16'b10111_111111_10101;
        tomato_soup[11][30] = 16'b10111_111111_10101;
        tomato_soup[11][31] = 16'b10111_111111_10101;
        tomato_soup[12][0] = 16'b10111_111111_10101;
        tomato_soup[12][1] = 16'b10111_111111_10101;
        tomato_soup[12][2] = 16'b10111_111111_10101;
        tomato_soup[12][3] = 16'b11001_101000_01100;
        tomato_soup[12][4] = 16'b11001_101001_01101;
        tomato_soup[12][5] = 16'b11011_101111_10001;
        tomato_soup[12][6] = 16'b11010_101011_01110;
        tomato_soup[12][7] = 16'b11000_010111_00100;
        tomato_soup[12][8] = 16'b10111_001011_00001;
        tomato_soup[12][9] = 16'b10110_001011_00001;
        tomato_soup[12][10] = 16'b10111_001011_00001;
        tomato_soup[12][11] = 16'b10111_001100_00001;
        tomato_soup[12][12] = 16'b10111_001100_00001;
        tomato_soup[12][13] = 16'b10111_001100_00001;
        tomato_soup[12][14] = 16'b11000_001110_00001;
        tomato_soup[12][15] = 16'b11001_001111_00001;
        tomato_soup[12][16] = 16'b11001_001110_00001;
        tomato_soup[12][17] = 16'b11000_001101_00001;
        tomato_soup[12][18] = 16'b11001_001111_00001;
        tomato_soup[12][19] = 16'b11000_001101_00001;
        tomato_soup[12][20] = 16'b11000_001101_00001;
        tomato_soup[12][21] = 16'b11000_001110_00001;
        tomato_soup[12][22] = 16'b10111_001100_00001;
        tomato_soup[12][23] = 16'b11000_010110_00100;
        tomato_soup[12][24] = 16'b11010_101010_01110;
        tomato_soup[12][25] = 16'b11011_110001_10010;
        tomato_soup[12][26] = 16'b11001_101001_01101;
        tomato_soup[12][27] = 16'b11001_101001_01101;
        tomato_soup[12][28] = 16'b10111_111111_10101;
        tomato_soup[12][29] = 16'b10111_111111_10101;
        tomato_soup[12][30] = 16'b10111_111111_10101;
        tomato_soup[12][31] = 16'b10111_111111_10101;
        tomato_soup[13][0] = 16'b10111_111111_10101;
        tomato_soup[13][1] = 16'b10111_111111_10101;
        tomato_soup[13][2] = 16'b10111_111111_10101;
        tomato_soup[13][3] = 16'b11001_101001_01101;
        tomato_soup[13][4] = 16'b11010_101101_01111;
        tomato_soup[13][5] = 16'b11001_011111_01000;
        tomato_soup[13][6] = 16'b10111_001100_00001;
        tomato_soup[13][7] = 16'b10111_001011_00001;
        tomato_soup[13][8] = 16'b10111_001100_00001;
        tomato_soup[13][9] = 16'b10111_001011_00001;
        tomato_soup[13][10] = 16'b11000_001110_00001;
        tomato_soup[13][11] = 16'b11000_001110_00001;
        tomato_soup[13][12] = 16'b11000_001110_00001;
        tomato_soup[13][13] = 16'b11000_001110_00001;
        tomato_soup[13][14] = 16'b11000_001110_00001;
        tomato_soup[13][15] = 16'b11001_001110_00001;
        tomato_soup[13][16] = 16'b11001_001111_00001;
        tomato_soup[13][17] = 16'b11001_001111_00001;
        tomato_soup[13][18] = 16'b11001_001111_00010;
        tomato_soup[13][19] = 16'b11000_001110_00001;
        tomato_soup[13][20] = 16'b11000_001110_00001;
        tomato_soup[13][21] = 16'b11000_001110_00001;
        tomato_soup[13][22] = 16'b11001_001110_00001;
        tomato_soup[13][23] = 16'b11000_001110_00001;
        tomato_soup[13][24] = 16'b11000_001101_00001;
        tomato_soup[13][25] = 16'b11001_100011_01010;
        tomato_soup[13][26] = 16'b11100_110001_10011;
        tomato_soup[13][27] = 16'b11001_101010_01101;
        tomato_soup[13][28] = 16'b11001_101001_01101;
        tomato_soup[13][29] = 16'b10111_111111_10101;
        tomato_soup[13][30] = 16'b10111_111111_10101;
        tomato_soup[13][31] = 16'b10111_111111_10101;
        tomato_soup[14][0] = 16'b10111_111111_10101;
        tomato_soup[14][1] = 16'b10111_111111_10101;
        tomato_soup[14][2] = 16'b11010_101110_10000;
        tomato_soup[14][3] = 16'b11011_101111_10001;
        tomato_soup[14][4] = 16'b11001_100010_01001;
        tomato_soup[14][5] = 16'b10111_001011_00001;
        tomato_soup[14][6] = 16'b10111_001100_00001;
        tomato_soup[14][7] = 16'b10111_001100_00001;
        tomato_soup[14][8] = 16'b11000_001110_00001;
        tomato_soup[14][9] = 16'b11001_001111_00010;
        tomato_soup[14][10] = 16'b11000_001101_00001;
        tomato_soup[14][11] = 16'b11001_001111_00010;
        tomato_soup[14][12] = 16'b11001_001111_00001;
        tomato_soup[14][13] = 16'b11000_001101_00001;
        tomato_soup[14][14] = 16'b11000_001110_00001;
        tomato_soup[14][15] = 16'b11000_001101_00001;
        tomato_soup[14][16] = 16'b10111_001100_00001;
        tomato_soup[14][17] = 16'b11000_001101_00001;
        tomato_soup[14][18] = 16'b10111_001100_00001;
        tomato_soup[14][19] = 16'b10111_001100_00001;
        tomato_soup[14][20] = 16'b10111_001100_00001;
        tomato_soup[14][21] = 16'b10111_001100_00001;
        tomato_soup[14][22] = 16'b11001_001110_00001;
        tomato_soup[14][23] = 16'b11001_001110_00010;
        tomato_soup[14][24] = 16'b11000_001110_00001;
        tomato_soup[14][25] = 16'b11000_001110_00001;
        tomato_soup[14][26] = 16'b11000_011011_00110;
        tomato_soup[14][27] = 16'b11011_110000_10010;
        tomato_soup[14][28] = 16'b11001_101001_01101;
        tomato_soup[14][29] = 16'b10111_111111_10101;
        tomato_soup[14][30] = 16'b10111_111111_10101;
        tomato_soup[14][31] = 16'b10111_111111_10101;
        tomato_soup[15][0] = 16'b10111_111111_10101;
        tomato_soup[15][1] = 16'b10111_111111_10101;
        tomato_soup[15][2] = 16'b11100_110010_10011;
        tomato_soup[15][3] = 16'b11100_110001_10011;
        tomato_soup[15][4] = 16'b10111_001100_00001;
        tomato_soup[15][5] = 16'b10111_001011_00001;
        tomato_soup[15][6] = 16'b10111_001100_00001;
        tomato_soup[15][7] = 16'b11000_001101_00001;
        tomato_soup[15][8] = 16'b11001_001110_00001;
        tomato_soup[15][9] = 16'b11010_010000_00010;
        tomato_soup[15][10] = 16'b11001_001110_00001;
        tomato_soup[15][11] = 16'b11000_001100_00001;
        tomato_soup[15][12] = 16'b11000_001110_00001;
        tomato_soup[15][13] = 16'b10111_001101_00001;
        tomato_soup[15][14] = 16'b11000_001101_00001;
        tomato_soup[15][15] = 16'b11000_001101_00001;
        tomato_soup[15][16] = 16'b11001_001110_00001;
        tomato_soup[15][17] = 16'b11001_001111_00001;
        tomato_soup[15][18] = 16'b11001_001110_00001;
        tomato_soup[15][19] = 16'b11000_001101_00001;
        tomato_soup[15][20] = 16'b10111_001100_00001;
        tomato_soup[15][21] = 16'b10111_001100_00001;
        tomato_soup[15][22] = 16'b10111_001100_00001;
        tomato_soup[15][23] = 16'b11000_001110_00001;
        tomato_soup[15][24] = 16'b11000_001110_00001;
        tomato_soup[15][25] = 16'b11001_001111_00001;
        tomato_soup[15][26] = 16'b10111_001011_00001;
        tomato_soup[15][27] = 16'b11001_100101_01011;
        tomato_soup[15][28] = 16'b11011_101110_10000;
        tomato_soup[15][29] = 16'b10111_111111_10101;
        tomato_soup[15][30] = 16'b10111_111111_10101;
        tomato_soup[15][31] = 16'b10111_111111_10101;
        tomato_soup[16][0] = 16'b10111_111111_10101;
        tomato_soup[16][1] = 16'b10111_111111_10101;
        tomato_soup[16][2] = 16'b11011_110001_10011;
        tomato_soup[16][3] = 16'b11011_110000_10010;
        tomato_soup[16][4] = 16'b10111_001011_00001;
        tomato_soup[16][5] = 16'b10111_001011_00001;
        tomato_soup[16][6] = 16'b10111_001100_00001;
        tomato_soup[16][7] = 16'b11001_001111_00010;
        tomato_soup[16][8] = 16'b11001_001111_00010;
        tomato_soup[16][9] = 16'b11001_001111_00010;
        tomato_soup[16][10] = 16'b11000_001101_00001;
        tomato_soup[16][11] = 16'b11000_001110_00001;
        tomato_soup[16][12] = 16'b11001_001111_00010;
        tomato_soup[16][13] = 16'b11000_001101_00001;
        tomato_soup[16][14] = 16'b11001_001111_00010;
        tomato_soup[16][15] = 16'b11001_001111_00001;
        tomato_soup[16][16] = 16'b11001_001111_00001;
        tomato_soup[16][17] = 16'b11001_001111_00010;
        tomato_soup[16][18] = 16'b11001_001111_00010;
        tomato_soup[16][19] = 16'b11000_001101_00001;
        tomato_soup[16][20] = 16'b10111_001100_00001;
        tomato_soup[16][21] = 16'b01100_011010_00011;
        tomato_soup[16][22] = 16'b01100_011010_00011;
        tomato_soup[16][23] = 16'b10111_001100_00001;
        tomato_soup[16][24] = 16'b11000_001101_00001;
        tomato_soup[16][25] = 16'b11001_001111_00010;
        tomato_soup[16][26] = 16'b10111_001011_00001;
        tomato_soup[16][27] = 16'b10111_010010_00011;
        tomato_soup[16][28] = 16'b11011_110000_10010;
        tomato_soup[16][29] = 16'b10111_111111_10101;
        tomato_soup[16][30] = 16'b10111_111111_10101;
        tomato_soup[16][31] = 16'b10111_111111_10101;
        tomato_soup[17][0] = 16'b10111_111111_10101;
        tomato_soup[17][1] = 16'b10111_111111_10101;
        tomato_soup[17][2] = 16'b11100_110010_10100;
        tomato_soup[17][3] = 16'b11010_101100_01111;
        tomato_soup[17][4] = 16'b10111_001110_00010;
        tomato_soup[17][5] = 16'b10111_001011_00001;
        tomato_soup[17][6] = 16'b10111_001100_00001;
        tomato_soup[17][7] = 16'b10111_001100_00001;
        tomato_soup[17][8] = 16'b11001_001111_00010;
        tomato_soup[17][9] = 16'b11001_001111_00010;
        tomato_soup[17][10] = 16'b11000_001101_00001;
        tomato_soup[17][11] = 16'b11000_001101_00001;
        tomato_soup[17][12] = 16'b11001_001111_00010;
        tomato_soup[17][13] = 16'b11000_001101_00001;
        tomato_soup[17][14] = 16'b11001_001111_00001;
        tomato_soup[17][15] = 16'b11001_001111_00010;
        tomato_soup[17][16] = 16'b11001_001111_00010;
        tomato_soup[17][17] = 16'b11000_001110_00001;
        tomato_soup[17][18] = 16'b11000_001110_00001;
        tomato_soup[17][19] = 16'b01100_011010_00011;
        tomato_soup[17][20] = 16'b01100_011001_00011;
        tomato_soup[17][21] = 16'b01100_011010_00011;
        tomato_soup[17][22] = 16'b01011_011001_00011;
        tomato_soup[17][23] = 16'b01011_010111_00010;
        tomato_soup[17][24] = 16'b10111_001100_00001;
        tomato_soup[17][25] = 16'b11001_010000_00010;
        tomato_soup[17][26] = 16'b10111_001011_00001;
        tomato_soup[17][27] = 16'b10111_010101_00100;
        tomato_soup[17][28] = 16'b11100_110010_10011;
        tomato_soup[17][29] = 16'b10111_111111_10101;
        tomato_soup[17][30] = 16'b10111_111111_10101;
        tomato_soup[17][31] = 16'b10111_111111_10101;
        tomato_soup[18][0] = 16'b10111_111111_10101;
        tomato_soup[18][1] = 16'b10111_111111_10101;
        tomato_soup[18][2] = 16'b11100_110010_10100;
        tomato_soup[18][3] = 16'b11010_101011_01110;
        tomato_soup[18][4] = 16'b11000_011100_00110;
        tomato_soup[18][5] = 16'b10111_001100_00001;
        tomato_soup[18][6] = 16'b10111_001011_00001;
        tomato_soup[18][7] = 16'b10111_001100_00001;
        tomato_soup[18][8] = 16'b11001_001111_00010;
        tomato_soup[18][9] = 16'b11001_001111_00001;
        tomato_soup[18][10] = 16'b11001_001111_00010;
        tomato_soup[18][11] = 16'b11000_001101_00001;
        tomato_soup[18][12] = 16'b11000_001101_00001;
        tomato_soup[18][13] = 16'b10111_001100_00001;
        tomato_soup[18][14] = 16'b11000_001101_00001;
        tomato_soup[18][15] = 16'b11000_001101_00001;
        tomato_soup[18][16] = 16'b11001_001110_00001;
        tomato_soup[18][17] = 16'b11000_001101_00001;
        tomato_soup[18][18] = 16'b01100_011010_00011;
        tomato_soup[18][19] = 16'b01100_011010_00011;
        tomato_soup[18][20] = 16'b01011_011001_00011;
        tomato_soup[18][21] = 16'b01101_011101_00011;
        tomato_soup[18][22] = 16'b01101_011101_00011;
        tomato_soup[18][23] = 16'b01100_011010_00011;
        tomato_soup[18][24] = 16'b10111_001100_00001;
        tomato_soup[18][25] = 16'b11000_001101_00001;
        tomato_soup[18][26] = 16'b10111_001011_00001;
        tomato_soup[18][27] = 16'b11001_101001_01101;
        tomato_soup[18][28] = 16'b11100_110010_10100;
        tomato_soup[18][29] = 16'b10111_111111_10101;
        tomato_soup[18][30] = 16'b10111_111111_10101;
        tomato_soup[18][31] = 16'b10111_111111_10101;
        tomato_soup[19][0] = 16'b10111_111111_10101;
        tomato_soup[19][1] = 16'b10111_111111_10101;
        tomato_soup[19][2] = 16'b10111_111111_10101;
        tomato_soup[19][3] = 16'b11011_101110_10000;
        tomato_soup[19][4] = 16'b11001_101001_01101;
        tomato_soup[19][5] = 16'b10111_011000_00101;
        tomato_soup[19][6] = 16'b10111_001100_00001;
        tomato_soup[19][7] = 16'b10111_001011_00001;
        tomato_soup[19][8] = 16'b11000_001110_00010;
        tomato_soup[19][9] = 16'b11001_001110_00001;
        tomato_soup[19][10] = 16'b11001_001111_00010;
        tomato_soup[19][11] = 16'b11000_001110_00001;
        tomato_soup[19][12] = 16'b11000_001110_00001;
        tomato_soup[19][13] = 16'b11000_001101_00001;
        tomato_soup[19][14] = 16'b11000_001101_00001;
        tomato_soup[19][15] = 16'b11000_001101_00001;
        tomato_soup[19][16] = 16'b11000_001101_00001;
        tomato_soup[19][17] = 16'b11000_001101_00001;
        tomato_soup[19][18] = 16'b01100_011010_00011;
        tomato_soup[19][19] = 16'b01100_011001_00011;
        tomato_soup[19][20] = 16'b01011_011001_00010;
        tomato_soup[19][21] = 16'b01010_010110_00010;
        tomato_soup[19][22] = 16'b01010_010101_00010;
        tomato_soup[19][23] = 16'b10111_001011_00001;
        tomato_soup[19][24] = 16'b10111_001100_00001;
        tomato_soup[19][25] = 16'b10111_001101_00001;
        tomato_soup[19][26] = 16'b11000_100000_01000;
        tomato_soup[19][27] = 16'b11010_101100_01111;
        tomato_soup[19][28] = 16'b11100_110011_10100;
        tomato_soup[19][29] = 16'b10111_111111_10101;
        tomato_soup[19][30] = 16'b10111_111111_10101;
        tomato_soup[19][31] = 16'b10111_111111_10101;
        tomato_soup[20][0] = 16'b10111_111111_10101;
        tomato_soup[20][1] = 16'b10111_111111_10101;
        tomato_soup[20][2] = 16'b10111_111111_10101;
        tomato_soup[20][3] = 16'b11010_101100_01111;
        tomato_soup[20][4] = 16'b11010_101011_01110;
        tomato_soup[20][5] = 16'b11001_101010_01110;
        tomato_soup[20][6] = 16'b11000_011110_00111;
        tomato_soup[20][7] = 16'b10111_001100_00001;
        tomato_soup[20][8] = 16'b10110_001011_00001;
        tomato_soup[20][9] = 16'b10111_001011_00001;
        tomato_soup[20][10] = 16'b11001_001111_00010;
        tomato_soup[20][11] = 16'b11001_001111_00010;
        tomato_soup[20][12] = 16'b11000_001110_00001;
        tomato_soup[20][13] = 16'b11000_001101_00001;
        tomato_soup[20][14] = 16'b11000_001110_00001;
        tomato_soup[20][15] = 16'b11001_001111_00001;
        tomato_soup[20][16] = 16'b11001_001111_00010;
        tomato_soup[20][17] = 16'b11001_001111_00001;
        tomato_soup[20][18] = 16'b11000_001110_00001;
        tomato_soup[20][19] = 16'b01100_011011_00011;
        tomato_soup[20][20] = 16'b01100_011010_00011;
        tomato_soup[20][21] = 16'b10111_001011_00001;
        tomato_soup[20][22] = 16'b10111_001011_00001;
        tomato_soup[20][23] = 16'b10111_001100_00001;
        tomato_soup[20][24] = 16'b10111_001100_00001;
        tomato_soup[20][25] = 16'b11001_100000_01000;
        tomato_soup[20][26] = 16'b11010_101010_01110;
        tomato_soup[20][27] = 16'b11011_101110_10001;
        tomato_soup[20][28] = 16'b11011_110000_10010;
        tomato_soup[20][29] = 16'b10111_111111_10101;
        tomato_soup[20][30] = 16'b10111_111111_10101;
        tomato_soup[20][31] = 16'b10111_111111_10101;
        tomato_soup[21][0] = 16'b10111_111111_10101;
        tomato_soup[21][1] = 16'b10111_111111_10101;
        tomato_soup[21][2] = 16'b10111_111111_10101;
        tomato_soup[21][3] = 16'b10111_111111_10101;
        tomato_soup[21][4] = 16'b11011_101110_10000;
        tomato_soup[21][5] = 16'b11001_101010_01110;
        tomato_soup[21][6] = 16'b11001_101001_01101;
        tomato_soup[21][7] = 16'b11001_101000_01100;
        tomato_soup[21][8] = 16'b10111_010100_00011;
        tomato_soup[21][9] = 16'b10111_001100_00001;
        tomato_soup[21][10] = 16'b10111_001100_00001;
        tomato_soup[21][11] = 16'b10111_001011_00000;
        tomato_soup[21][12] = 16'b10111_001011_00001;
        tomato_soup[21][13] = 16'b10111_001011_00000;
        tomato_soup[21][14] = 16'b10111_001100_00001;
        tomato_soup[21][15] = 16'b11001_001110_00001;
        tomato_soup[21][16] = 16'b11001_001111_00001;
        tomato_soup[21][17] = 16'b11001_001110_00001;
        tomato_soup[21][18] = 16'b11001_001110_00001;
        tomato_soup[21][19] = 16'b11000_001100_00001;
        tomato_soup[21][20] = 16'b10111_001100_00001;
        tomato_soup[21][21] = 16'b10111_001100_00001;
        tomato_soup[21][22] = 16'b10111_001100_00001;
        tomato_soup[21][23] = 16'b11000_010110_00100;
        tomato_soup[21][24] = 16'b11001_101001_01101;
        tomato_soup[21][25] = 16'b11001_101001_01101;
        tomato_soup[21][26] = 16'b11010_101011_01110;
        tomato_soup[21][27] = 16'b11011_110000_10010;
        tomato_soup[21][28] = 16'b10111_111111_10101;
        tomato_soup[21][29] = 16'b10111_111111_10101;
        tomato_soup[21][30] = 16'b10111_111111_10101;
        tomato_soup[21][31] = 16'b10111_111111_10101;
        tomato_soup[22][0] = 16'b10111_111111_10101;
        tomato_soup[22][1] = 16'b10111_111111_10101;
        tomato_soup[22][2] = 16'b10111_111111_10101;
        tomato_soup[22][3] = 16'b10111_111111_10101;
        tomato_soup[22][4] = 16'b10111_111111_10101;
        tomato_soup[22][5] = 16'b11011_110001_10010;
        tomato_soup[22][6] = 16'b11001_101010_01101;
        tomato_soup[22][7] = 16'b11001_101001_01101;
        tomato_soup[22][8] = 16'b11001_101001_01101;
        tomato_soup[22][9] = 16'b11001_101000_01100;
        tomato_soup[22][10] = 16'b11001_101000_01100;
        tomato_soup[22][11] = 16'b11000_010100_00011;
        tomato_soup[22][12] = 16'b10111_001100_00001;
        tomato_soup[22][13] = 16'b10111_001011_00001;
        tomato_soup[22][14] = 16'b10111_001100_00001;
        tomato_soup[22][15] = 16'b10111_001100_00001;
        tomato_soup[22][16] = 16'b10111_001100_00001;
        tomato_soup[22][17] = 16'b11001_001110_00001;
        tomato_soup[22][18] = 16'b11000_001110_00001;
        tomato_soup[22][19] = 16'b11000_001101_00001;
        tomato_soup[22][20] = 16'b11000_010110_00100;
        tomato_soup[22][21] = 16'b11001_101000_01100;
        tomato_soup[22][22] = 16'b11001_101000_01100;
        tomato_soup[22][23] = 16'b11001_101001_01101;
        tomato_soup[22][24] = 16'b11001_101001_01101;
        tomato_soup[22][25] = 16'b11001_101010_01110;
        tomato_soup[22][26] = 16'b11011_101111_10001;
        tomato_soup[22][27] = 16'b10111_111111_10101;
        tomato_soup[22][28] = 16'b10111_111111_10101;
        tomato_soup[22][29] = 16'b10111_111111_10101;
        tomato_soup[22][30] = 16'b10111_111111_10101;
        tomato_soup[22][31] = 16'b10111_111111_10101;
        tomato_soup[23][0] = 16'b10111_111111_10101;
        tomato_soup[23][1] = 16'b10111_111111_10101;
        tomato_soup[23][2] = 16'b10111_111111_10101;
        tomato_soup[23][3] = 16'b10111_111111_10101;
        tomato_soup[23][4] = 16'b10111_111111_10101;
        tomato_soup[23][5] = 16'b10111_111111_10101;
        tomato_soup[23][6] = 16'b11011_101110_10000;
        tomato_soup[23][7] = 16'b11010_101110_10000;
        tomato_soup[23][8] = 16'b11001_101001_01101;
        tomato_soup[23][9] = 16'b11001_101001_01101;
        tomato_soup[23][10] = 16'b11001_101010_01101;
        tomato_soup[23][11] = 16'b11001_101001_01101;
        tomato_soup[23][12] = 16'b11001_101000_01101;
        tomato_soup[23][13] = 16'b11001_101000_01100;
        tomato_soup[23][14] = 16'b11001_101001_01101;
        tomato_soup[23][15] = 16'b11001_101001_01101;
        tomato_soup[23][16] = 16'b11001_101000_01100;
        tomato_soup[23][17] = 16'b11001_101001_01101;
        tomato_soup[23][18] = 16'b11001_101001_01101;
        tomato_soup[23][19] = 16'b11001_101000_01100;
        tomato_soup[23][20] = 16'b11001_101000_01101;
        tomato_soup[23][21] = 16'b11001_101001_01101;
        tomato_soup[23][22] = 16'b11001_101001_01101;
        tomato_soup[23][23] = 16'b11010_101101_01111;
        tomato_soup[23][24] = 16'b11011_101111_10001;
        tomato_soup[23][25] = 16'b11011_101110_10000;
        tomato_soup[23][26] = 16'b10111_111111_10101;
        tomato_soup[23][27] = 16'b10111_111111_10101;
        tomato_soup[23][28] = 16'b10111_111111_10101;
        tomato_soup[23][29] = 16'b10111_111111_10101;
        tomato_soup[23][30] = 16'b10111_111111_10101;
        tomato_soup[23][31] = 16'b10111_111111_10101;
        tomato_soup[24][0] = 16'b10111_111111_10101;
        tomato_soup[24][1] = 16'b10111_111111_10101;
        tomato_soup[24][2] = 16'b10111_111111_10101;
        tomato_soup[24][3] = 16'b10111_111111_10101;
        tomato_soup[24][4] = 16'b10111_111111_10101;
        tomato_soup[24][5] = 16'b10111_111111_10101;
        tomato_soup[24][6] = 16'b10111_111111_10101;
        tomato_soup[24][7] = 16'b11011_110000_10010;
        tomato_soup[24][8] = 16'b11011_110001_10011;
        tomato_soup[24][9] = 16'b11011_110000_10010;
        tomato_soup[24][10] = 16'b11011_110000_10010;
        tomato_soup[24][11] = 16'b11001_101001_01101;
        tomato_soup[24][12] = 16'b11001_101001_01101;
        tomato_soup[24][13] = 16'b11001_101000_01100;
        tomato_soup[24][14] = 16'b11001_101000_01100;
        tomato_soup[24][15] = 16'b11001_101000_01100;
        tomato_soup[24][16] = 16'b11001_101000_01100;
        tomato_soup[24][17] = 16'b11001_101001_01101;
        tomato_soup[24][18] = 16'b11001_101001_01101;
        tomato_soup[24][19] = 16'b11001_101000_01100;
        tomato_soup[24][20] = 16'b11001_101001_01101;
        tomato_soup[24][21] = 16'b11010_101110_10000;
        tomato_soup[24][22] = 16'b11011_110001_10010;
        tomato_soup[24][23] = 16'b11011_110001_10011;
        tomato_soup[24][24] = 16'b11011_110000_10010;
        tomato_soup[24][25] = 16'b10111_111111_10101;
        tomato_soup[24][26] = 16'b10111_111111_10101;
        tomato_soup[24][27] = 16'b10111_111111_10101;
        tomato_soup[24][28] = 16'b10111_111111_10101;
        tomato_soup[24][29] = 16'b10111_111111_10101;
        tomato_soup[24][30] = 16'b10111_111111_10101;
        tomato_soup[24][31] = 16'b10111_111111_10101;
        tomato_soup[25][0] = 16'b10110_111111_10100;
        tomato_soup[25][1] = 16'b10111_111111_10101;
        tomato_soup[25][2] = 16'b10111_111111_10101;
        tomato_soup[25][3] = 16'b10111_111111_10101;
        tomato_soup[25][4] = 16'b10111_111111_10101;
        tomato_soup[25][5] = 16'b10111_111111_10101;
        tomato_soup[25][6] = 16'b10111_111111_10101;
        tomato_soup[25][7] = 16'b10111_111111_10101;
        tomato_soup[25][8] = 16'b10111_111111_10101;
        tomato_soup[25][9] = 16'b10111_111111_10101;
        tomato_soup[25][10] = 16'b11100_110010_10011;
        tomato_soup[25][11] = 16'b11100_110010_10011;
        tomato_soup[25][12] = 16'b11011_110001_10010;
        tomato_soup[25][13] = 16'b11100_110010_10011;
        tomato_soup[25][14] = 16'b11011_110001_10010;
        tomato_soup[25][15] = 16'b11011_110001_10010;
        tomato_soup[25][16] = 16'b11011_110001_10010;
        tomato_soup[25][17] = 16'b11011_110001_10010;
        tomato_soup[25][18] = 16'b11011_110001_10010;
        tomato_soup[25][19] = 16'b11011_101110_10001;
        tomato_soup[25][20] = 16'b11011_110000_10010;
        tomato_soup[25][21] = 16'b11011_110001_10010;
        tomato_soup[25][22] = 16'b10111_111111_10101;
        tomato_soup[25][23] = 16'b10111_111111_10101;
        tomato_soup[25][24] = 16'b10111_111111_10101;
        tomato_soup[25][25] = 16'b10111_111111_10101;
        tomato_soup[25][26] = 16'b10111_111111_10101;
        tomato_soup[25][27] = 16'b10111_111111_10101;
        tomato_soup[25][28] = 16'b10111_111111_10101;
        tomato_soup[25][29] = 16'b10111_111111_10101;
        tomato_soup[25][30] = 16'b10111_111111_10101;
        tomato_soup[25][31] = 16'b10111_111111_10101;
        tomato_soup[26][0] = 16'b10111_111111_10101;
        tomato_soup[26][1] = 16'b10111_111111_10101;
        tomato_soup[26][2] = 16'b10110_111111_10100;
        tomato_soup[26][3] = 16'b10111_111111_10101;
        tomato_soup[26][4] = 16'b10111_111111_10101;
        tomato_soup[26][5] = 16'b10111_111111_10101;
        tomato_soup[26][6] = 16'b10111_111111_10101;
        tomato_soup[26][7] = 16'b10111_111111_10101;
        tomato_soup[26][8] = 16'b10111_111111_10101;
        tomato_soup[26][9] = 16'b10111_111111_10101;
        tomato_soup[26][10] = 16'b10111_111111_10101;
        tomato_soup[26][11] = 16'b10111_111111_10101;
        tomato_soup[26][12] = 16'b10111_111111_10101;
        tomato_soup[26][13] = 16'b10111_111111_10101;
        tomato_soup[26][14] = 16'b10111_111111_10101;
        tomato_soup[26][15] = 16'b10111_111111_10101;
        tomato_soup[26][16] = 16'b10111_111111_10101;
        tomato_soup[26][17] = 16'b10111_111111_10101;
        tomato_soup[26][18] = 16'b10111_111111_10101;
        tomato_soup[26][19] = 16'b10111_111111_10101;
        tomato_soup[26][20] = 16'b10111_111111_10101;
        tomato_soup[26][21] = 16'b10111_111111_10101;
        tomato_soup[26][22] = 16'b10111_111111_10101;
        tomato_soup[26][23] = 16'b10111_111111_10101;
        tomato_soup[26][24] = 16'b10111_111111_10101;
        tomato_soup[26][25] = 16'b10111_111111_10101;
        tomato_soup[26][26] = 16'b10111_111111_10101;
        tomato_soup[26][27] = 16'b10111_111111_10101;
        tomato_soup[26][28] = 16'b10111_111111_10101;
        tomato_soup[26][29] = 16'b10111_111111_10101;
        tomato_soup[26][30] = 16'b10111_111111_10101;
        tomato_soup[26][31] = 16'b10111_111111_10101;
        tomato_soup[27][0] = 16'b10111_111111_10101;
        tomato_soup[27][1] = 16'b10111_111111_10101;
        tomato_soup[27][2] = 16'b10111_111111_10101;
        tomato_soup[27][3] = 16'b10110_111111_10100;
        tomato_soup[27][4] = 16'b10111_111111_10101;
        tomato_soup[27][5] = 16'b10111_111111_10101;
        tomato_soup[27][6] = 16'b10111_111111_10101;
        tomato_soup[27][7] = 16'b10111_111111_10101;
        tomato_soup[27][8] = 16'b10111_111111_10101;
        tomato_soup[27][9] = 16'b10111_111111_10101;
        tomato_soup[27][10] = 16'b10111_111111_10101;
        tomato_soup[27][11] = 16'b10111_111111_10101;
        tomato_soup[27][12] = 16'b10111_111111_10101;
        tomato_soup[27][13] = 16'b10111_111111_10101;
        tomato_soup[27][14] = 16'b10111_111111_10101;
        tomato_soup[27][15] = 16'b10111_111111_10101;
        tomato_soup[27][16] = 16'b10111_111111_10101;
        tomato_soup[27][17] = 16'b10111_111111_10101;
        tomato_soup[27][18] = 16'b10111_111111_10101;
        tomato_soup[27][19] = 16'b10111_111111_10101;
        tomato_soup[27][20] = 16'b10111_111111_10101;
        tomato_soup[27][21] = 16'b10111_111111_10101;
        tomato_soup[27][22] = 16'b10111_111111_10101;
        tomato_soup[27][23] = 16'b10111_111111_10101;
        tomato_soup[27][24] = 16'b10111_111111_10101;
        tomato_soup[27][25] = 16'b10111_111111_10101;
        tomato_soup[27][26] = 16'b10111_111111_10101;
        tomato_soup[27][27] = 16'b10111_111111_10101;
        tomato_soup[27][28] = 16'b10111_111111_10101;
        tomato_soup[27][29] = 16'b10111_111111_10101;
        tomato_soup[27][30] = 16'b10111_111111_10101;
        tomato_soup[27][31] = 16'b10111_111111_10101;
        tomato_soup[28][0] = 16'b10111_111111_10101;
        tomato_soup[28][1] = 16'b10111_111111_10101;
        tomato_soup[28][2] = 16'b10111_111111_10101;
        tomato_soup[28][3] = 16'b10110_111111_10100;
        tomato_soup[28][4] = 16'b10111_111111_10101;
        tomato_soup[28][5] = 16'b10111_111111_10101;
        tomato_soup[28][6] = 16'b10111_111111_10101;
        tomato_soup[28][7] = 16'b10111_111111_10101;
        tomato_soup[28][8] = 16'b10111_111111_10101;
        tomato_soup[28][9] = 16'b10111_111111_10101;
        tomato_soup[28][10] = 16'b10111_111111_10101;
        tomato_soup[28][11] = 16'b10111_111111_10101;
        tomato_soup[28][12] = 16'b10111_111111_10101;
        tomato_soup[28][13] = 16'b10111_111111_10101;
        tomato_soup[28][14] = 16'b10111_111111_10101;
        tomato_soup[28][15] = 16'b10111_111111_10101;
        tomato_soup[28][16] = 16'b10111_111111_10101;
        tomato_soup[28][17] = 16'b10111_111111_10101;
        tomato_soup[28][18] = 16'b10111_111111_10101;
        tomato_soup[28][19] = 16'b10111_111111_10101;
        tomato_soup[28][20] = 16'b10111_111111_10101;
        tomato_soup[28][21] = 16'b10111_111111_10101;
        tomato_soup[28][22] = 16'b10111_111111_10101;
        tomato_soup[28][23] = 16'b10111_111111_10101;
        tomato_soup[28][24] = 16'b10111_111111_10101;
        tomato_soup[28][25] = 16'b10111_111111_10101;
        tomato_soup[28][26] = 16'b10111_111111_10101;
        tomato_soup[28][27] = 16'b10111_111111_10101;
        tomato_soup[28][28] = 16'b10111_111111_10101;
        tomato_soup[28][29] = 16'b10111_111111_10101;
        tomato_soup[28][30] = 16'b10111_111111_10101;
        tomato_soup[28][31] = 16'b10111_111111_10101;
        tomato_soup[29][0] = 16'b10111_111111_10101;
        tomato_soup[29][1] = 16'b10111_111111_10101;
        tomato_soup[29][2] = 16'b10111_111111_10101;
        tomato_soup[29][3] = 16'b10111_111111_10101;
        tomato_soup[29][4] = 16'b10111_111111_10101;
        tomato_soup[29][5] = 16'b10111_111111_10101;
        tomato_soup[29][6] = 16'b10111_111111_10101;
        tomato_soup[29][7] = 16'b10111_111111_10101;
        tomato_soup[29][8] = 16'b10111_111111_10101;
        tomato_soup[29][9] = 16'b10111_111111_10101;
        tomato_soup[29][10] = 16'b10111_111111_10101;
        tomato_soup[29][11] = 16'b10111_111111_10101;
        tomato_soup[29][12] = 16'b10111_111111_10101;
        tomato_soup[29][13] = 16'b10111_111111_10101;
        tomato_soup[29][14] = 16'b10111_111111_10101;
        tomato_soup[29][15] = 16'b10111_111111_10101;
        tomato_soup[29][16] = 16'b10111_111111_10101;
        tomato_soup[29][17] = 16'b10111_111111_10101;
        tomato_soup[29][18] = 16'b10111_111111_10101;
        tomato_soup[29][19] = 16'b10111_111111_10101;
        tomato_soup[29][20] = 16'b10111_111111_10101;
        tomato_soup[29][21] = 16'b10111_111111_10101;
        tomato_soup[29][22] = 16'b10111_111111_10101;
        tomato_soup[29][23] = 16'b10111_111111_10101;
        tomato_soup[29][24] = 16'b10111_111111_10101;
        tomato_soup[29][25] = 16'b10111_111111_10101;
        tomato_soup[29][26] = 16'b10111_111111_10101;
        tomato_soup[29][27] = 16'b10111_111111_10101;
        tomato_soup[29][28] = 16'b10111_111111_10101;
        tomato_soup[29][29] = 16'b10111_111111_10101;
        tomato_soup[29][30] = 16'b10111_111111_10101;
        tomato_soup[29][31] = 16'b10111_111111_10101;
        tomato_soup[30][0] = 16'b10111_111111_10101;
        tomato_soup[30][1] = 16'b10111_111111_10101;
        tomato_soup[30][2] = 16'b10111_111111_10101;
        tomato_soup[30][3] = 16'b10111_111111_10101;
        tomato_soup[30][4] = 16'b10111_111111_10101;
        tomato_soup[30][5] = 16'b10111_111111_10101;
        tomato_soup[30][6] = 16'b10111_111111_10101;
        tomato_soup[30][7] = 16'b10111_111111_10101;
        tomato_soup[30][8] = 16'b10111_111111_10101;
        tomato_soup[30][9] = 16'b10111_111111_10101;
        tomato_soup[30][10] = 16'b10111_111111_10101;
        tomato_soup[30][11] = 16'b10111_111111_10101;
        tomato_soup[30][12] = 16'b10111_111111_10101;
        tomato_soup[30][13] = 16'b10111_111111_10101;
        tomato_soup[30][14] = 16'b10111_111111_10101;
        tomato_soup[30][15] = 16'b10111_111111_10101;
        tomato_soup[30][16] = 16'b10111_111111_10101;
        tomato_soup[30][17] = 16'b10111_111111_10101;
        tomato_soup[30][18] = 16'b10111_111111_10101;
        tomato_soup[30][19] = 16'b10111_111111_10101;
        tomato_soup[30][20] = 16'b10111_111111_10101;
        tomato_soup[30][21] = 16'b10111_111111_10101;
        tomato_soup[30][22] = 16'b10111_111111_10101;
        tomato_soup[30][23] = 16'b10111_111111_10101;
        tomato_soup[30][24] = 16'b10111_111111_10101;
        tomato_soup[30][25] = 16'b10111_111111_10101;
        tomato_soup[30][26] = 16'b10111_111111_10101;
        tomato_soup[30][27] = 16'b10111_111111_10101;
        tomato_soup[30][28] = 16'b10111_111111_10101;
        tomato_soup[30][29] = 16'b10111_111111_10101;
        tomato_soup[30][30] = 16'b10111_111111_10101;
        tomato_soup[30][31] = 16'b10111_111111_10101;
        tomato_soup[31][0] = 16'b10111_111111_10101;
        tomato_soup[31][1] = 16'b10111_111111_10101;
        tomato_soup[31][2] = 16'b10111_111111_10101;
        tomato_soup[31][3] = 16'b10111_111111_10101;
        tomato_soup[31][4] = 16'b10111_111111_10101;
        tomato_soup[31][5] = 16'b10111_111111_10101;
        tomato_soup[31][6] = 16'b10111_111111_10101;
        tomato_soup[31][7] = 16'b10111_111111_10101;
        tomato_soup[31][8] = 16'b10111_111111_10101;
        tomato_soup[31][9] = 16'b10111_111111_10101;
        tomato_soup[31][10] = 16'b10111_111111_10101;
        tomato_soup[31][11] = 16'b10111_111111_10101;
        tomato_soup[31][12] = 16'b10111_111111_10101;
        tomato_soup[31][13] = 16'b10111_111111_10101;
        tomato_soup[31][14] = 16'b10111_111111_10101;
        tomato_soup[31][15] = 16'b10111_111111_10101;
        tomato_soup[31][16] = 16'b10111_111111_10101;
        tomato_soup[31][17] = 16'b10111_111111_10101;
        tomato_soup[31][18] = 16'b10111_111111_10101;
        tomato_soup[31][19] = 16'b10111_111111_10101;
        tomato_soup[31][20] = 16'b10111_111111_10101;
        tomato_soup[31][21] = 16'b10111_111111_10101;
        tomato_soup[31][22] = 16'b10111_111111_10101;
        tomato_soup[31][23] = 16'b10111_111111_10101;
        tomato_soup[31][24] = 16'b10111_111111_10101;
        tomato_soup[31][25] = 16'b10111_111111_10101;
        tomato_soup[31][26] = 16'b10111_111111_10101;
        tomato_soup[31][27] = 16'b10111_111111_10101;
        tomato_soup[31][28] = 16'b10111_111111_10101;
        tomato_soup[31][29] = 16'b10111_111111_10101;
        tomato_soup[31][30] = 16'b10111_111111_10101;
        tomato_soup[31][31] = 16'b10111_111111_10101;



        tomato_rice[0][0] = 16'b11110_110000_11110;
        tomato_rice[0][1] = 16'b11110_110000_11110;
        tomato_rice[0][2] = 16'b11110_110000_11110;
        tomato_rice[0][3] = 16'b11110_110000_11110;
        tomato_rice[0][4] = 16'b11110_110000_11110;
        tomato_rice[0][5] = 16'b11110_110000_11110;
        tomato_rice[0][6] = 16'b11110_110000_11110;
        tomato_rice[0][7] = 16'b11110_110000_11110;
        tomato_rice[0][8] = 16'b11110_110000_11110;
        tomato_rice[0][9] = 16'b11110_110000_11110;
        tomato_rice[0][10] = 16'b11110_110000_11110;
        tomato_rice[0][11] = 16'b11110_110000_11110;
        tomato_rice[0][12] = 16'b11110_110000_11110;
        tomato_rice[0][13] = 16'b11110_110000_11110;
        tomato_rice[0][14] = 16'b11110_110000_11110;
        tomato_rice[0][15] = 16'b11110_110000_11110;
        tomato_rice[0][16] = 16'b11110_110000_11110;
        tomato_rice[0][17] = 16'b11110_110000_11110;
        tomato_rice[0][18] = 16'b11110_110000_11110;
        tomato_rice[0][19] = 16'b11110_110000_11110;
        tomato_rice[0][20] = 16'b11110_110000_11110;
        tomato_rice[0][21] = 16'b11110_110000_11110;
        tomato_rice[0][22] = 16'b11110_110000_11110;
        tomato_rice[0][23] = 16'b11110_110000_11110;
        tomato_rice[0][24] = 16'b11110_110000_11110;
        tomato_rice[0][25] = 16'b11110_110000_11110;
        tomato_rice[0][26] = 16'b11110_110000_11110;
        tomato_rice[0][27] = 16'b11110_110000_11110;
        tomato_rice[0][28] = 16'b11110_110000_11110;
        tomato_rice[0][29] = 16'b11110_110000_11110;
        tomato_rice[0][30] = 16'b11110_110000_11110;
        tomato_rice[0][31] = 16'b11110_110000_11110;
        tomato_rice[1][0] = 16'b11110_110000_11110;
        tomato_rice[1][1] = 16'b11110_110000_11110;
        tomato_rice[1][2] = 16'b11110_110000_11110;
        tomato_rice[1][3] = 16'b11110_110000_11110;
        tomato_rice[1][4] = 16'b11110_110000_11110;
        tomato_rice[1][5] = 16'b11110_110000_11110;
        tomato_rice[1][6] = 16'b11110_110000_11110;
        tomato_rice[1][7] = 16'b11110_110000_11110;
        tomato_rice[1][8] = 16'b11110_110000_11110;
        tomato_rice[1][9] = 16'b11110_110000_11110;
        tomato_rice[1][10] = 16'b11110_110000_11110;
        tomato_rice[1][11] = 16'b11110_110000_11110;
        tomato_rice[1][12] = 16'b11110_110000_11110;
        tomato_rice[1][13] = 16'b11110_110000_11110;
        tomato_rice[1][14] = 16'b11110_110000_11110;
        tomato_rice[1][15] = 16'b11110_110000_11110;
        tomato_rice[1][16] = 16'b11110_110000_11110;
        tomato_rice[1][17] = 16'b11110_110000_11110;
        tomato_rice[1][18] = 16'b11110_110000_11110;
        tomato_rice[1][19] = 16'b11110_110000_11110;
        tomato_rice[1][20] = 16'b11110_110000_11110;
        tomato_rice[1][21] = 16'b11110_110000_11110;
        tomato_rice[1][22] = 16'b11110_110000_11110;
        tomato_rice[1][23] = 16'b11110_110000_11110;
        tomato_rice[1][24] = 16'b11110_110000_11110;
        tomato_rice[1][25] = 16'b11110_110000_11110;
        tomato_rice[1][26] = 16'b11110_110000_11110;
        tomato_rice[1][27] = 16'b11110_110000_11110;
        tomato_rice[1][28] = 16'b11110_110000_11110;
        tomato_rice[1][29] = 16'b11110_110000_11110;
        tomato_rice[1][30] = 16'b11110_110000_11110;
        tomato_rice[1][31] = 16'b11110_110000_11110;
        tomato_rice[2][0] = 16'b11110_110000_11110;
        tomato_rice[2][1] = 16'b11110_110000_11110;
        tomato_rice[2][2] = 16'b11110_110000_11110;
        tomato_rice[2][3] = 16'b11110_110000_11110;
        tomato_rice[2][4] = 16'b11110_110000_11110;
        tomato_rice[2][5] = 16'b11110_110000_11110;
        tomato_rice[2][6] = 16'b11110_110000_11110;
        tomato_rice[2][7] = 16'b11110_110000_11110;
        tomato_rice[2][8] = 16'b11110_110000_11110;
        tomato_rice[2][9] = 16'b11110_110000_11110;
        tomato_rice[2][10] = 16'b11110_110000_11110;
        tomato_rice[2][11] = 16'b11110_110000_11110;
        tomato_rice[2][12] = 16'b11110_110000_11110;
        tomato_rice[2][13] = 16'b11110_110000_11110;
        tomato_rice[2][14] = 16'b11110_110000_11110;
        tomato_rice[2][15] = 16'b11110_110000_11110;
        tomato_rice[2][16] = 16'b11110_110000_11110;
        tomato_rice[2][17] = 16'b11110_110000_11110;
        tomato_rice[2][18] = 16'b11110_110000_11110;
        tomato_rice[2][19] = 16'b11110_110000_11110;
        tomato_rice[2][20] = 16'b11110_110000_11110;
        tomato_rice[2][21] = 16'b11110_110000_11110;
        tomato_rice[2][22] = 16'b11110_110000_11110;
        tomato_rice[2][23] = 16'b11110_110000_11110;
        tomato_rice[2][24] = 16'b11110_110000_11110;
        tomato_rice[2][25] = 16'b11110_110000_11110;
        tomato_rice[2][26] = 16'b11110_110000_11110;
        tomato_rice[2][27] = 16'b11110_110000_11110;
        tomato_rice[2][28] = 16'b11110_110000_11110;
        tomato_rice[2][29] = 16'b11110_110000_11110;
        tomato_rice[2][30] = 16'b11110_110000_11110;
        tomato_rice[2][31] = 16'b11110_110000_11110;
        tomato_rice[3][0] = 16'b11110_110000_11110;
        tomato_rice[3][1] = 16'b11110_110000_11110;
        tomato_rice[3][2] = 16'b11110_110000_11110;
        tomato_rice[3][3] = 16'b11110_110000_11110;
        tomato_rice[3][4] = 16'b11110_110000_11110;
        tomato_rice[3][5] = 16'b11110_110000_11110;
        tomato_rice[3][6] = 16'b11110_110000_11110;
        tomato_rice[3][7] = 16'b11110_110000_11110;
        tomato_rice[3][8] = 16'b11110_110000_11110;
        tomato_rice[3][9] = 16'b11110_110000_11110;
        tomato_rice[3][10] = 16'b11110_110000_11110;
        tomato_rice[3][11] = 16'b11110_110000_11110;
        tomato_rice[3][12] = 16'b11110_110000_11110;
        tomato_rice[3][13] = 16'b11110_110000_11110;
        tomato_rice[3][14] = 16'b11110_110000_11110;
        tomato_rice[3][15] = 16'b11110_110000_11110;
        tomato_rice[3][16] = 16'b11110_110000_11110;
        tomato_rice[3][17] = 16'b11110_110000_11110;
        tomato_rice[3][18] = 16'b11110_110000_11110;
        tomato_rice[3][19] = 16'b11110_110000_11110;
        tomato_rice[3][20] = 16'b11110_110000_11110;
        tomato_rice[3][21] = 16'b11110_110000_11110;
        tomato_rice[3][22] = 16'b11110_110000_11110;
        tomato_rice[3][23] = 16'b11110_110000_11110;
        tomato_rice[3][24] = 16'b11110_110000_11110;
        tomato_rice[3][25] = 16'b11110_110000_11110;
        tomato_rice[3][26] = 16'b11110_110000_11110;
        tomato_rice[3][27] = 16'b11110_110000_11110;
        tomato_rice[3][28] = 16'b11110_110000_11110;
        tomato_rice[3][29] = 16'b11110_110000_11110;
        tomato_rice[3][30] = 16'b11110_110000_11110;
        tomato_rice[3][31] = 16'b11110_110000_11110;
        tomato_rice[4][0] = 16'b11110_110000_11110;
        tomato_rice[4][1] = 16'b11110_110000_11110;
        tomato_rice[4][2] = 16'b11110_110000_11110;
        tomato_rice[4][3] = 16'b11110_110000_11110;
        tomato_rice[4][4] = 16'b11110_110000_11110;
        tomato_rice[4][5] = 16'b11110_110000_11110;
        tomato_rice[4][6] = 16'b11110_110000_11110;
        tomato_rice[4][7] = 16'b11110_110000_11110;
        tomato_rice[4][8] = 16'b11110_110000_11110;
        tomato_rice[4][9] = 16'b11110_110000_11110;
        tomato_rice[4][10] = 16'b11110_110000_11110;
        tomato_rice[4][11] = 16'b11110_110000_11110;
        tomato_rice[4][12] = 16'b11110_110000_11110;
        tomato_rice[4][13] = 16'b11110_110000_11110;
        tomato_rice[4][14] = 16'b11110_110000_11110;
        tomato_rice[4][15] = 16'b11110_110000_11110;
        tomato_rice[4][16] = 16'b11110_110000_11110;
        tomato_rice[4][17] = 16'b11110_110000_11110;
        tomato_rice[4][18] = 16'b11110_110000_11110;
        tomato_rice[4][19] = 16'b11110_110000_11110;
        tomato_rice[4][20] = 16'b11110_110000_11110;
        tomato_rice[4][21] = 16'b11110_110000_11110;
        tomato_rice[4][22] = 16'b11110_110000_11110;
        tomato_rice[4][23] = 16'b11110_110000_11110;
        tomato_rice[4][24] = 16'b11110_110000_11110;
        tomato_rice[4][25] = 16'b11110_110000_11110;
        tomato_rice[4][26] = 16'b11110_110000_11110;
        tomato_rice[4][27] = 16'b11110_110000_11110;
        tomato_rice[4][28] = 16'b11110_110000_11110;
        tomato_rice[4][29] = 16'b11110_110000_11110;
        tomato_rice[4][30] = 16'b11110_110000_11110;
        tomato_rice[4][31] = 16'b11110_110000_11110;
        tomato_rice[5][0] = 16'b11110_110000_11110;
        tomato_rice[5][1] = 16'b11110_110000_11110;
        tomato_rice[5][2] = 16'b11110_110000_11110;
        tomato_rice[5][3] = 16'b11110_110000_11110;
        tomato_rice[5][4] = 16'b11110_110000_11110;
        tomato_rice[5][5] = 16'b11110_110000_11110;
        tomato_rice[5][6] = 16'b11110_110000_11110;
        tomato_rice[5][7] = 16'b11110_110000_11110;
        tomato_rice[5][8] = 16'b11110_110000_11110;
        tomato_rice[5][9] = 16'b11110_110000_11110;
        tomato_rice[5][10] = 16'b11001_101001_01101;
        tomato_rice[5][11] = 16'b11001_101000_01100;
        tomato_rice[5][12] = 16'b11001_101001_01100;
        tomato_rice[5][13] = 16'b11001_101001_01100;
        tomato_rice[5][14] = 16'b11001_101001_01101;
        tomato_rice[5][15] = 16'b11010_101101_01110;
        tomato_rice[5][16] = 16'b11010_101011_01110;
        tomato_rice[5][17] = 16'b11010_101010_01101;
        tomato_rice[5][18] = 16'b11010_101010_01101;
        tomato_rice[5][19] = 16'b11001_101010_01101;
        tomato_rice[5][20] = 16'b11001_101010_01101;
        tomato_rice[5][21] = 16'b11001_101010_01101;
        tomato_rice[5][22] = 16'b11110_110000_11110;
        tomato_rice[5][23] = 16'b11110_110000_11110;
        tomato_rice[5][24] = 16'b11110_110000_11110;
        tomato_rice[5][25] = 16'b11110_110000_11110;
        tomato_rice[5][26] = 16'b11110_110000_11110;
        tomato_rice[5][27] = 16'b11110_110000_11110;
        tomato_rice[5][28] = 16'b11110_110000_11110;
        tomato_rice[5][29] = 16'b11110_110000_11110;
        tomato_rice[5][30] = 16'b11110_110000_11110;
        tomato_rice[5][31] = 16'b11110_110000_11110;
        tomato_rice[6][0] = 16'b11110_110000_11110;
        tomato_rice[6][1] = 16'b11110_110000_11110;
        tomato_rice[6][2] = 16'b11110_110000_11110;
        tomato_rice[6][3] = 16'b11110_110000_11110;
        tomato_rice[6][4] = 16'b11110_110000_11110;
        tomato_rice[6][5] = 16'b11110_110000_11110;
        tomato_rice[6][6] = 16'b11110_110000_11110;
        tomato_rice[6][7] = 16'b11001_101001_01101;
        tomato_rice[6][8] = 16'b11001_101000_01100;
        tomato_rice[6][9] = 16'b11011_101110_01111;
        tomato_rice[6][10] = 16'b11011_110000_10000;
        tomato_rice[6][11] = 16'b11011_110000_10000;
        tomato_rice[6][12] = 16'b11011_101111_10000;
        tomato_rice[6][13] = 16'b11100_110000_10001;
        tomato_rice[6][14] = 16'b11011_101110_10000;
        tomato_rice[6][15] = 16'b11011_101101_01111;
        tomato_rice[6][16] = 16'b11011_101111_10000;
        tomato_rice[6][17] = 16'b11011_101110_10000;
        tomato_rice[6][18] = 16'b11011_101111_10000;
        tomato_rice[6][19] = 16'b11011_101111_10000;
        tomato_rice[6][20] = 16'b11011_101111_10000;
        tomato_rice[6][21] = 16'b11011_101101_01111;
        tomato_rice[6][22] = 16'b11010_101010_01101;
        tomato_rice[6][23] = 16'b11010_101011_01110;
        tomato_rice[6][24] = 16'b11001_101001_01101;
        tomato_rice[6][25] = 16'b11110_110000_11110;
        tomato_rice[6][26] = 16'b11110_110000_11110;
        tomato_rice[6][27] = 16'b11110_110000_11110;
        tomato_rice[6][28] = 16'b11110_110000_11110;
        tomato_rice[6][29] = 16'b11110_110000_11110;
        tomato_rice[6][30] = 16'b11110_110000_11110;
        tomato_rice[6][31] = 16'b11110_110000_11110;
        tomato_rice[7][0] = 16'b11110_110000_11110;
        tomato_rice[7][1] = 16'b11110_110000_11110;
        tomato_rice[7][2] = 16'b11110_110000_11110;
        tomato_rice[7][3] = 16'b11110_110000_11110;
        tomato_rice[7][4] = 16'b11110_110000_11110;
        tomato_rice[7][5] = 16'b11001_101000_01100;
        tomato_rice[7][6] = 16'b11001_101001_01100;
        tomato_rice[7][7] = 16'b11011_101111_10000;
        tomato_rice[7][8] = 16'b11011_101111_10000;
        tomato_rice[7][9] = 16'b11011_101110_10000;
        tomato_rice[7][10] = 16'b11011_101110_01111;
        tomato_rice[7][11] = 16'b11011_110000_10000;
        tomato_rice[7][12] = 16'b11011_101110_10000;
        tomato_rice[7][13] = 16'b11011_101110_10000;
        tomato_rice[7][14] = 16'b11011_101110_10000;
        tomato_rice[7][15] = 16'b11011_101101_01111;
        tomato_rice[7][16] = 16'b11011_101101_01111;
        tomato_rice[7][17] = 16'b11011_101110_01111;
        tomato_rice[7][18] = 16'b11011_101101_01111;
        tomato_rice[7][19] = 16'b11010_101101_01111;
        tomato_rice[7][20] = 16'b11011_101110_01111;
        tomato_rice[7][21] = 16'b11011_101111_10000;
        tomato_rice[7][22] = 16'b11011_101110_01111;
        tomato_rice[7][23] = 16'b11011_101111_10000;
        tomato_rice[7][24] = 16'b11011_101111_10000;
        tomato_rice[7][25] = 16'b11001_101001_01101;
        tomato_rice[7][26] = 16'b11001_101001_01100;
        tomato_rice[7][27] = 16'b11110_110000_11110;
        tomato_rice[7][28] = 16'b11110_110000_11110;
        tomato_rice[7][29] = 16'b11110_110000_11110;
        tomato_rice[7][30] = 16'b11110_110000_11110;
        tomato_rice[7][31] = 16'b11110_110000_11110;
        tomato_rice[8][0] = 16'b11110_110000_11110;
        tomato_rice[8][1] = 16'b11110_110000_11110;
        tomato_rice[8][2] = 16'b11110_110000_11110;
        tomato_rice[8][3] = 16'b11110_110000_11110;
        tomato_rice[8][4] = 16'b11001_100111_01011;
        tomato_rice[8][5] = 16'b11011_101110_01111;
        tomato_rice[8][6] = 16'b11011_110000_10000;
        tomato_rice[8][7] = 16'b11100_110000_10001;
        tomato_rice[8][8] = 16'b11011_101110_01111;
        tomato_rice[8][9] = 16'b11011_101101_01111;
        tomato_rice[8][10] = 16'b11011_110000_10000;
        tomato_rice[8][11] = 16'b11011_101111_10000;
        tomato_rice[8][12] = 16'b11010_101011_01110;
        tomato_rice[8][13] = 16'b11001_101000_01100;
        tomato_rice[8][14] = 16'b11010_101001_01100;
        tomato_rice[8][15] = 16'b11010_101001_01100;
        tomato_rice[8][16] = 16'b11001_101001_01100;
        tomato_rice[8][17] = 16'b11001_100110_01010;
        tomato_rice[8][18] = 16'b11000_100101_01010;
        tomato_rice[8][19] = 16'b11010_101011_01110;
        tomato_rice[8][20] = 16'b11011_101111_10000;
        tomato_rice[8][21] = 16'b11011_101110_01111;
        tomato_rice[8][22] = 16'b11011_101110_01111;
        tomato_rice[8][23] = 16'b11011_101111_10000;
        tomato_rice[8][24] = 16'b11011_110000_10000;
        tomato_rice[8][25] = 16'b11100_110000_10000;
        tomato_rice[8][26] = 16'b11011_101110_10000;
        tomato_rice[8][27] = 16'b11001_101001_01101;
        tomato_rice[8][28] = 16'b11110_110000_11110;
        tomato_rice[8][29] = 16'b11110_110000_11110;
        tomato_rice[8][30] = 16'b11110_110000_11110;
        tomato_rice[8][31] = 16'b11110_110000_11110;
        tomato_rice[9][0] = 16'b11110_110000_11110;
        tomato_rice[9][1] = 16'b11110_110000_11110;
        tomato_rice[9][2] = 16'b11110_110000_11110;
        tomato_rice[9][3] = 16'b11001_101001_01101;
        tomato_rice[9][4] = 16'b11011_101110_10000;
        tomato_rice[9][5] = 16'b11011_101110_10000;
        tomato_rice[9][6] = 16'b11011_101111_10000;
        tomato_rice[9][7] = 16'b11011_110000_10001;
        tomato_rice[9][8] = 16'b11011_101111_10000;
        tomato_rice[9][9] = 16'b11010_101010_01101;
        tomato_rice[9][10] = 16'b11010_101010_01101;
        tomato_rice[9][11] = 16'b11010_101010_01101;
        tomato_rice[9][12] = 16'b11001_100001_01001;
        tomato_rice[9][13] = 16'b11001_011011_00101;
        tomato_rice[9][14] = 16'b11001_010111_00100;
        tomato_rice[9][15] = 16'b11000_001111_00001;
        tomato_rice[9][16] = 16'b11000_001111_00001;
        tomato_rice[9][17] = 16'b11001_010110_00011;
        tomato_rice[9][18] = 16'b11001_011000_00100;
        tomato_rice[9][19] = 16'b11001_100101_01011;
        tomato_rice[9][20] = 16'b11001_101001_01101;
        tomato_rice[9][21] = 16'b11010_101010_01101;
        tomato_rice[9][22] = 16'b11010_101010_01101;
        tomato_rice[9][23] = 16'b11011_101110_01111;
        tomato_rice[9][24] = 16'b11011_101111_10000;
        tomato_rice[9][25] = 16'b11011_101111_10000;
        tomato_rice[9][26] = 16'b11011_101111_10000;
        tomato_rice[9][27] = 16'b11100_110001_10001;
        tomato_rice[9][28] = 16'b11001_101010_01101;
        tomato_rice[9][29] = 16'b11110_110000_11110;
        tomato_rice[9][30] = 16'b11110_110000_11110;
        tomato_rice[9][31] = 16'b11110_110000_11110;
        tomato_rice[10][0] = 16'b11110_110000_11110;
        tomato_rice[10][1] = 16'b11110_110000_11110;
        tomato_rice[10][2] = 16'b11110_110000_11110;
        tomato_rice[10][3] = 16'b11011_101111_10000;
        tomato_rice[10][4] = 16'b11011_101111_10000;
        tomato_rice[10][5] = 16'b11011_101111_10000;
        tomato_rice[10][6] = 16'b11011_101110_01111;
        tomato_rice[10][7] = 16'b11010_101010_01101;
        tomato_rice[10][8] = 16'b11010_101001_01100;
        tomato_rice[10][9] = 16'b11010_100000_01000;
        tomato_rice[10][10] = 16'b11010_011011_00110;
        tomato_rice[10][11] = 16'b11001_010001_00010;
        tomato_rice[10][12] = 16'b11001_010001_00001;
        tomato_rice[10][13] = 16'b11010_010011_00010;
        tomato_rice[10][14] = 16'b11001_010010_00010;
        tomato_rice[10][15] = 16'b11000_010000_00001;
        tomato_rice[10][16] = 16'b11001_010011_00010;
        tomato_rice[10][17] = 16'b11001_010011_00010;
        tomato_rice[10][18] = 16'b11010_010101_00011;
        tomato_rice[10][19] = 16'b11010_010100_00010;
        tomato_rice[10][20] = 16'b11001_010010_00010;
        tomato_rice[10][21] = 16'b11001_010001_00001;
        tomato_rice[10][22] = 16'b11010_011101_00110;
        tomato_rice[10][23] = 16'b11010_101010_01101;
        tomato_rice[10][24] = 16'b11001_101000_01100;
        tomato_rice[10][25] = 16'b11011_101111_10000;
        tomato_rice[10][26] = 16'b11100_110000_10001;
        tomato_rice[10][27] = 16'b11011_101111_10000;
        tomato_rice[10][28] = 16'b11011_101111_10000;
        tomato_rice[10][29] = 16'b11110_110000_11110;
        tomato_rice[10][30] = 16'b11110_110000_11110;
        tomato_rice[10][31] = 16'b11110_110000_11110;
        tomato_rice[11][0] = 16'b11110_110000_11110;
        tomato_rice[11][1] = 16'b11110_110000_11110;
        tomato_rice[11][2] = 16'b11010_101011_01110;
        tomato_rice[11][3] = 16'b11011_101111_10000;
        tomato_rice[11][4] = 16'b11100_110000_10001;
        tomato_rice[11][5] = 16'b11011_110000_10001;
        tomato_rice[11][6] = 16'b11010_101010_01101;
        tomato_rice[11][7] = 16'b11010_011101_00110;
        tomato_rice[11][8] = 16'b11001_010001_00001;
        tomato_rice[11][9] = 16'b11000_010000_00001;
        tomato_rice[11][10] = 16'b11000_001111_00001;
        tomato_rice[11][11] = 16'b11010_010100_00010;
        tomato_rice[11][12] = 16'b11010_010100_00010;
        tomato_rice[11][13] = 16'b11001_010010_00010;
        tomato_rice[11][14] = 16'b11011_010110_00011;
        tomato_rice[11][15] = 16'b11010_010101_00011;
        tomato_rice[11][16] = 16'b11010_010101_00011;
        tomato_rice[11][17] = 16'b11001_010010_00010;
        tomato_rice[11][18] = 16'b11001_010010_00010;
        tomato_rice[11][19] = 16'b11001_010010_00010;
        tomato_rice[11][20] = 16'b11010_010011_00010;
        tomato_rice[11][21] = 16'b11001_010010_00001;
        tomato_rice[11][22] = 16'b11001_010010_00010;
        tomato_rice[11][23] = 16'b11001_010001_00010;
        tomato_rice[11][24] = 16'b11001_011110_00111;
        tomato_rice[11][25] = 16'b11010_101001_01100;
        tomato_rice[11][26] = 16'b11011_101110_10000;
        tomato_rice[11][27] = 16'b11011_101110_01111;
        tomato_rice[11][28] = 16'b11011_101110_01111;
        tomato_rice[11][29] = 16'b11011_101101_01111;
        tomato_rice[11][30] = 16'b11110_110000_11110;
        tomato_rice[11][31] = 16'b11110_110000_11110;
        tomato_rice[12][0] = 16'b11110_110000_11110;
        tomato_rice[12][1] = 16'b11110_110000_11110;
        tomato_rice[12][2] = 16'b11011_110000_10000;
        tomato_rice[12][3] = 16'b11011_101110_10000;
        tomato_rice[12][4] = 16'b11011_101111_10000;
        tomato_rice[12][5] = 16'b11010_101010_01101;
        tomato_rice[12][6] = 16'b11001_011011_00101;
        tomato_rice[12][7] = 16'b11000_010000_00001;
        tomato_rice[12][8] = 16'b11001_010000_00001;
        tomato_rice[12][9] = 16'b11010_010011_00010;
        tomato_rice[12][10] = 16'b11010_010011_00010;
        tomato_rice[12][11] = 16'b11000_001111_00001;
        tomato_rice[12][12] = 16'b11010_010011_00010;
        tomato_rice[12][13] = 16'b11010_010011_00010;
        tomato_rice[12][14] = 16'b11001_010010_00010;
        tomato_rice[12][15] = 16'b11010_010101_00010;
        tomato_rice[12][16] = 16'b11010_010010_00010;
        tomato_rice[12][17] = 16'b11010_010011_00010;
        tomato_rice[12][18] = 16'b11011_010101_00011;
        tomato_rice[12][19] = 16'b11010_010101_00010;
        tomato_rice[12][20] = 16'b11001_010001_00001;
        tomato_rice[12][21] = 16'b11001_010001_00010;
        tomato_rice[12][22] = 16'b11001_010010_00010;
        tomato_rice[12][23] = 16'b11010_010011_00010;
        tomato_rice[12][24] = 16'b11001_010000_00001;
        tomato_rice[12][25] = 16'b11001_011001_00101;
        tomato_rice[12][26] = 16'b11010_101001_01101;
        tomato_rice[12][27] = 16'b11011_101111_10000;
        tomato_rice[12][28] = 16'b11011_101110_01111;
        tomato_rice[12][29] = 16'b11011_101111_10000;
        tomato_rice[12][30] = 16'b11110_110000_11110;
        tomato_rice[12][31] = 16'b11110_110000_11110;
        tomato_rice[13][0] = 16'b11110_110000_11110;
        tomato_rice[13][1] = 16'b11110_110000_11110;
        tomato_rice[13][2] = 16'b11011_101111_10000;
        tomato_rice[13][3] = 16'b11011_110000_10001;
        tomato_rice[13][4] = 16'b11100_110000_10001;
        tomato_rice[13][5] = 16'b11001_101001_01100;
        tomato_rice[13][6] = 16'b11000_001111_00001;
        tomato_rice[13][7] = 16'b11010_010011_00010;
        tomato_rice[13][8] = 16'b11010_010011_00010;
        tomato_rice[13][9] = 16'b11001_010000_00001;
        tomato_rice[13][10] = 16'b11010_010011_00010;
        tomato_rice[13][11] = 16'b11010_010011_00010;
        tomato_rice[13][12] = 16'b11001_010000_00001;
        tomato_rice[13][13] = 16'b11010_010101_00011;
        tomato_rice[13][14] = 16'b11010_010101_00010;
        tomato_rice[13][15] = 16'b11010_010010_00010;
        tomato_rice[13][16] = 16'b11011_010111_00011;
        tomato_rice[13][17] = 16'b11011_010101_00011;
        tomato_rice[13][18] = 16'b11011_010110_00011;
        tomato_rice[13][19] = 16'b11010_010010_00010;
        tomato_rice[13][20] = 16'b11010_010100_00010;
        tomato_rice[13][21] = 16'b11010_010010_00010;
        tomato_rice[13][22] = 16'b11010_010010_00010;
        tomato_rice[13][23] = 16'b11011_011000_00100;
        tomato_rice[13][24] = 16'b11010_010011_00010;
        tomato_rice[13][25] = 16'b11001_010001_00010;
        tomato_rice[13][26] = 16'b11001_101000_01100;
        tomato_rice[13][27] = 16'b11100_110000_10000;
        tomato_rice[13][28] = 16'b11011_101111_10000;
        tomato_rice[13][29] = 16'b11011_110000_10000;
        tomato_rice[13][30] = 16'b11110_110000_11110;
        tomato_rice[13][31] = 16'b11110_110000_11110;
        tomato_rice[14][0] = 16'b11110_110000_11110;
        tomato_rice[14][1] = 16'b11110_110000_11110;
        tomato_rice[14][2] = 16'b11011_101111_10000;
        tomato_rice[14][3] = 16'b11011_101111_10000;
        tomato_rice[14][4] = 16'b11011_101111_10000;
        tomato_rice[14][5] = 16'b11001_101000_01100;
        tomato_rice[14][6] = 16'b11001_010011_00010;
        tomato_rice[14][7] = 16'b11001_010010_00010;
        tomato_rice[14][8] = 16'b11001_010010_00010;
        tomato_rice[14][9] = 16'b11010_010011_00010;
        tomato_rice[14][10] = 16'b11010_010010_00010;
        tomato_rice[14][11] = 16'b11011_010111_00011;
        tomato_rice[14][12] = 16'b11010_010100_00010;
        tomato_rice[14][13] = 16'b11011_010101_00011;
        tomato_rice[14][14] = 16'b11011_011000_00011;
        tomato_rice[14][15] = 16'b11011_010101_00011;
        tomato_rice[14][16] = 16'b11011_010101_00011;
        tomato_rice[14][17] = 16'b11010_010101_00010;
        tomato_rice[14][18] = 16'b11010_010010_00010;
        tomato_rice[14][19] = 16'b11010_010100_00010;
        tomato_rice[14][20] = 16'b11011_010101_00011;
        tomato_rice[14][21] = 16'b11011_010110_00011;
        tomato_rice[14][22] = 16'b11010_010100_00010;
        tomato_rice[14][23] = 16'b11010_010011_00010;
        tomato_rice[14][24] = 16'b11010_010011_00010;
        tomato_rice[14][25] = 16'b11010_010101_00011;
        tomato_rice[14][26] = 16'b11010_101010_01101;
        tomato_rice[14][27] = 16'b11011_101111_10000;
        tomato_rice[14][28] = 16'b11011_101101_01111;
        tomato_rice[14][29] = 16'b11100_110001_10001;
        tomato_rice[14][30] = 16'b11110_110000_11110;
        tomato_rice[14][31] = 16'b11110_110000_11110;
        tomato_rice[15][0] = 16'b11110_110000_11110;
        tomato_rice[15][1] = 16'b11110_110000_11110;
        tomato_rice[15][2] = 16'b11011_101111_10000;
        tomato_rice[15][3] = 16'b11011_101111_10000;
        tomato_rice[15][4] = 16'b11011_101111_10000;
        tomato_rice[15][5] = 16'b11010_101011_01110;
        tomato_rice[15][6] = 16'b11010_010111_00011;
        tomato_rice[15][7] = 16'b11001_010001_00001;
        tomato_rice[15][8] = 16'b11010_010010_00010;
        tomato_rice[15][9] = 16'b11100_011001_00100;
        tomato_rice[15][10] = 16'b11011_011000_00100;
        tomato_rice[15][11] = 16'b11010_010010_00010;
        tomato_rice[15][12] = 16'b11011_011000_00011;
        tomato_rice[15][13] = 16'b11010_010101_00010;
        tomato_rice[15][14] = 16'b11011_010110_00011;
        tomato_rice[15][15] = 16'b11010_010100_00010;
        tomato_rice[15][16] = 16'b11100_011010_00100;
        tomato_rice[15][17] = 16'b11100_011010_00100;
        tomato_rice[15][18] = 16'b11100_011001_00100;
        tomato_rice[15][19] = 16'b11011_010111_00011;
        tomato_rice[15][20] = 16'b11010_010011_00010;
        tomato_rice[15][21] = 16'b11010_010100_00010;
        tomato_rice[15][22] = 16'b11011_010111_00011;
        tomato_rice[15][23] = 16'b11011_011000_00100;
        tomato_rice[15][24] = 16'b11010_010011_00010;
        tomato_rice[15][25] = 16'b11010_010101_00010;
        tomato_rice[15][26] = 16'b11011_101110_01111;
        tomato_rice[15][27] = 16'b11011_101110_01111;
        tomato_rice[15][28] = 16'b11011_101101_01111;
        tomato_rice[15][29] = 16'b11011_101110_10000;
        tomato_rice[15][30] = 16'b11110_110000_11110;
        tomato_rice[15][31] = 16'b11110_110000_11110;
        tomato_rice[16][0] = 16'b11110_110000_11110;
        tomato_rice[16][1] = 16'b11110_110000_11110;
        tomato_rice[16][2] = 16'b11110_110000_11110;
        tomato_rice[16][3] = 16'b11011_101101_01111;
        tomato_rice[16][4] = 16'b11011_101110_01111;
        tomato_rice[16][5] = 16'b11011_101101_01111;
        tomato_rice[16][6] = 16'b11011_100011_01001;
        tomato_rice[16][7] = 16'b11010_010101_00011;
        tomato_rice[16][8] = 16'b11011_010101_00011;
        tomato_rice[16][9] = 16'b11010_010100_00010;
        tomato_rice[16][10] = 16'b11100_011001_00100;
        tomato_rice[16][11] = 16'b11011_010110_00011;
        tomato_rice[16][12] = 16'b11011_011000_00011;
        tomato_rice[16][13] = 16'b11011_011001_00100;
        tomato_rice[16][14] = 16'b11011_010110_00011;
        tomato_rice[16][15] = 16'b11011_010111_00011;
        tomato_rice[16][16] = 16'b11011_010101_00010;
        tomato_rice[16][17] = 16'b11011_011001_00100;
        tomato_rice[16][18] = 16'b11010_010101_00010;
        tomato_rice[16][19] = 16'b11011_010111_00011;
        tomato_rice[16][20] = 16'b11010_010100_00010;
        tomato_rice[16][21] = 16'b11010_010011_00010;
        tomato_rice[16][22] = 16'b11010_010101_00011;
        tomato_rice[16][23] = 16'b11011_010110_00011;
        tomato_rice[16][24] = 16'b11010_010101_00011;
        tomato_rice[16][25] = 16'b11011_100001_01000;
        tomato_rice[16][26] = 16'b11100_110000_10001;
        tomato_rice[16][27] = 16'b11011_101110_01111;
        tomato_rice[16][28] = 16'b11011_101110_10000;
        tomato_rice[16][29] = 16'b11110_110000_11110;
        tomato_rice[16][30] = 16'b11110_110000_11110;
        tomato_rice[16][31] = 16'b11110_110000_11110;
        tomato_rice[17][0] = 16'b11110_110000_11110;
        tomato_rice[17][1] = 16'b11110_110000_11110;
        tomato_rice[17][2] = 16'b11110_110000_11110;
        tomato_rice[17][3] = 16'b11110_110000_11110;
        tomato_rice[17][4] = 16'b11011_101101_01111;
        tomato_rice[17][5] = 16'b11010_101101_01111;
        tomato_rice[17][6] = 16'b11011_101110_01111;
        tomato_rice[17][7] = 16'b11001_010001_00010;
        tomato_rice[17][8] = 16'b11011_010101_00011;
        tomato_rice[17][9] = 16'b11011_010110_00011;
        tomato_rice[17][10] = 16'b11100_011001_00100;
        tomato_rice[17][11] = 16'b11011_010111_00011;
        tomato_rice[17][12] = 16'b11011_010101_00011;
        tomato_rice[17][13] = 16'b11011_011000_00100;
        tomato_rice[17][14] = 16'b11100_011110_00110;
        tomato_rice[17][15] = 16'b11011_011000_00100;
        tomato_rice[17][16] = 16'b11011_010110_00011;
        tomato_rice[17][17] = 16'b11011_010111_00011;
        tomato_rice[17][18] = 16'b11011_011001_00100;
        tomato_rice[17][19] = 16'b11011_010111_00011;
        tomato_rice[17][20] = 16'b11011_010111_00011;
        tomato_rice[17][21] = 16'b11011_011001_00100;
        tomato_rice[17][22] = 16'b11011_010111_00011;
        tomato_rice[17][23] = 16'b11001_010001_00001;
        tomato_rice[17][24] = 16'b11010_010101_00011;
        tomato_rice[17][25] = 16'b11011_101100_01110;
        tomato_rice[17][26] = 16'b11011_101110_01111;
        tomato_rice[17][27] = 16'b11011_110000_10000;
        tomato_rice[17][28] = 16'b11110_110000_11110;
        tomato_rice[17][29] = 16'b11110_110000_11110;
        tomato_rice[17][30] = 16'b11110_110000_11110;
        tomato_rice[17][31] = 16'b11110_110000_11110;
        tomato_rice[18][0] = 16'b11110_110000_11110;
        tomato_rice[18][1] = 16'b11110_110000_11110;
        tomato_rice[18][2] = 16'b11110_110000_11110;
        tomato_rice[18][3] = 16'b11110_110000_11110;
        tomato_rice[18][4] = 16'b11110_110000_11110;
        tomato_rice[18][5] = 16'b11011_101101_01111;
        tomato_rice[18][6] = 16'b11011_101101_01111;
        tomato_rice[18][7] = 16'b11010_010101_00011;
        tomato_rice[18][8] = 16'b11010_010011_00010;
        tomato_rice[18][9] = 16'b11011_010110_00011;
        tomato_rice[18][10] = 16'b11010_010011_00010;
        tomato_rice[18][11] = 16'b11011_010111_00011;
        tomato_rice[18][12] = 16'b11011_011000_00100;
        tomato_rice[18][13] = 16'b11011_011010_00100;
        tomato_rice[18][14] = 16'b11011_011001_00100;
        tomato_rice[18][15] = 16'b11011_010111_00011;
        tomato_rice[18][16] = 16'b11100_011010_00100;
        tomato_rice[18][17] = 16'b11011_010111_00011;
        tomato_rice[18][18] = 16'b11011_011001_00100;
        tomato_rice[18][19] = 16'b11100_011010_00100;
        tomato_rice[18][20] = 16'b11011_010110_00011;
        tomato_rice[18][21] = 16'b11010_010010_00010;
        tomato_rice[18][22] = 16'b11010_010101_00010;
        tomato_rice[18][23] = 16'b11011_010111_00011;
        tomato_rice[18][24] = 16'b11010_010101_00010;
        tomato_rice[18][25] = 16'b11011_101101_01110;
        tomato_rice[18][26] = 16'b11011_101110_01111;
        tomato_rice[18][27] = 16'b11110_110000_11110;
        tomato_rice[18][28] = 16'b11110_110000_11110;
        tomato_rice[18][29] = 16'b11110_110000_11110;
        tomato_rice[18][30] = 16'b11110_110000_11110;
        tomato_rice[18][31] = 16'b11110_110000_11110;
        tomato_rice[19][0] = 16'b11110_110000_11110;
        tomato_rice[19][1] = 16'b11110_110000_11110;
        tomato_rice[19][2] = 16'b11110_110000_11110;
        tomato_rice[19][3] = 16'b11110_110000_11110;
        tomato_rice[19][4] = 16'b11110_110000_11110;
        tomato_rice[19][5] = 16'b11110_110000_11110;
        tomato_rice[19][6] = 16'b11110_110000_11110;
        tomato_rice[19][7] = 16'b11100_100100_01010;
        tomato_rice[19][8] = 16'b11011_010101_00011;
        tomato_rice[19][9] = 16'b11011_010110_00011;
        tomato_rice[19][10] = 16'b11011_011000_00011;
        tomato_rice[19][11] = 16'b11011_011000_00100;
        tomato_rice[19][12] = 16'b11011_010100_00010;
        tomato_rice[19][13] = 16'b11011_011001_00100;
        tomato_rice[19][14] = 16'b11100_011111_00111;
        tomato_rice[19][15] = 16'b11011_011001_00100;
        tomato_rice[19][16] = 16'b11011_011001_00100;
        tomato_rice[19][17] = 16'b11011_011000_00100;
        tomato_rice[19][18] = 16'b11011_011000_00100;
        tomato_rice[19][19] = 16'b11011_010111_00011;
        tomato_rice[19][20] = 16'b11011_011000_00011;
        tomato_rice[19][21] = 16'b11010_010010_00010;
        tomato_rice[19][22] = 16'b11011_010101_00011;
        tomato_rice[19][23] = 16'b11011_010110_00011;
        tomato_rice[19][24] = 16'b11100_100100_01001;
        tomato_rice[19][25] = 16'b11110_110000_11110;
        tomato_rice[19][26] = 16'b11110_110000_11110;
        tomato_rice[19][27] = 16'b11110_110000_11110;
        tomato_rice[19][28] = 16'b11110_110000_11110;
        tomato_rice[19][29] = 16'b11110_110000_11110;
        tomato_rice[19][30] = 16'b11110_110000_11110;
        tomato_rice[19][31] = 16'b11110_110000_11110;
        tomato_rice[20][0] = 16'b11110_110000_11110;
        tomato_rice[20][1] = 16'b11110_110000_11110;
        tomato_rice[20][2] = 16'b11110_110000_11110;
        tomato_rice[20][3] = 16'b11110_110000_11110;
        tomato_rice[20][4] = 16'b11110_110000_11110;
        tomato_rice[20][5] = 16'b11110_110000_11110;
        tomato_rice[20][6] = 16'b11110_110000_11110;
        tomato_rice[20][7] = 16'b11110_110000_11110;
        tomato_rice[20][8] = 16'b11011_011000_00100;
        tomato_rice[20][9] = 16'b11011_010101_00010;
        tomato_rice[20][10] = 16'b11011_010111_00011;
        tomato_rice[20][11] = 16'b11011_011000_00011;
        tomato_rice[20][12] = 16'b11011_011001_00100;
        tomato_rice[20][13] = 16'b11011_011001_00100;
        tomato_rice[20][14] = 16'b11011_010110_00011;
        tomato_rice[20][15] = 16'b11011_011000_00011;
        tomato_rice[20][16] = 16'b11100_011100_00101;
        tomato_rice[20][17] = 16'b11011_011000_00100;
        tomato_rice[20][18] = 16'b11011_010110_00011;
        tomato_rice[20][19] = 16'b11100_011101_00101;
        tomato_rice[20][20] = 16'b11011_011000_00100;
        tomato_rice[20][21] = 16'b11011_010110_00011;
        tomato_rice[20][22] = 16'b11010_010010_00010;
        tomato_rice[20][23] = 16'b11011_010110_00011;
        tomato_rice[20][24] = 16'b11110_110000_11110;
        tomato_rice[20][25] = 16'b11110_110000_11110;
        tomato_rice[20][26] = 16'b11110_110000_11110;
        tomato_rice[20][27] = 16'b11110_110000_11110;
        tomato_rice[20][28] = 16'b11110_110000_11110;
        tomato_rice[20][29] = 16'b11110_110000_11110;
        tomato_rice[20][30] = 16'b11110_110000_11110;
        tomato_rice[20][31] = 16'b11110_110000_11110;
        tomato_rice[21][0] = 16'b11110_110000_11110;
        tomato_rice[21][1] = 16'b11110_110000_11110;
        tomato_rice[21][2] = 16'b11110_110000_11110;
        tomato_rice[21][3] = 16'b11110_110000_11110;
        tomato_rice[21][4] = 16'b11110_110000_11110;
        tomato_rice[21][5] = 16'b11110_110000_11110;
        tomato_rice[21][6] = 16'b11110_110000_11110;
        tomato_rice[21][7] = 16'b11110_110000_11110;
        tomato_rice[21][8] = 16'b11110_110000_11110;
        tomato_rice[21][9] = 16'b11011_011000_00100;
        tomato_rice[21][10] = 16'b11011_010110_00011;
        tomato_rice[21][11] = 16'b11100_011011_00101;
        tomato_rice[21][12] = 16'b11100_011010_00100;
        tomato_rice[21][13] = 16'b11010_010100_00010;
        tomato_rice[21][14] = 16'b11011_011000_00011;
        tomato_rice[21][15] = 16'b11100_011100_00101;
        tomato_rice[21][16] = 16'b11100_011101_00101;
        tomato_rice[21][17] = 16'b11011_010110_00011;
        tomato_rice[21][18] = 16'b11100_011010_00100;
        tomato_rice[21][19] = 16'b11011_010110_00011;
        tomato_rice[21][20] = 16'b11100_011001_00100;
        tomato_rice[21][21] = 16'b11100_011010_00100;
        tomato_rice[21][22] = 16'b11011_010111_00011;
        tomato_rice[21][23] = 16'b11110_110000_11110;
        tomato_rice[21][24] = 16'b11110_110000_11110;
        tomato_rice[21][25] = 16'b11110_110000_11110;
        tomato_rice[21][26] = 16'b11110_110000_11110;
        tomato_rice[21][27] = 16'b11110_110000_11110;
        tomato_rice[21][28] = 16'b11110_110000_11110;
        tomato_rice[21][29] = 16'b11110_110000_11110;
        tomato_rice[21][30] = 16'b11110_110000_11110;
        tomato_rice[21][31] = 16'b11110_110000_11110;
        tomato_rice[22][0] = 16'b11110_110000_11110;
        tomato_rice[22][1] = 16'b11110_110000_11110;
        tomato_rice[22][2] = 16'b11110_110000_11110;
        tomato_rice[22][3] = 16'b11110_110000_11110;
        tomato_rice[22][4] = 16'b11110_110000_11110;
        tomato_rice[22][5] = 16'b11110_110000_11110;
        tomato_rice[22][6] = 16'b11110_110000_11110;
        tomato_rice[22][7] = 16'b11110_110000_11110;
        tomato_rice[22][8] = 16'b11110_110000_11110;
        tomato_rice[22][9] = 16'b11110_110000_11110;
        tomato_rice[22][10] = 16'b11100_010111_00011;
        tomato_rice[22][11] = 16'b11011_010110_00011;
        tomato_rice[22][12] = 16'b11100_011011_00101;
        tomato_rice[22][13] = 16'b11100_011010_00100;
        tomato_rice[22][14] = 16'b11011_010110_00011;
        tomato_rice[22][15] = 16'b11011_011000_00011;
        tomato_rice[22][16] = 16'b11100_011001_00100;
        tomato_rice[22][17] = 16'b11100_011001_00100;
        tomato_rice[22][18] = 16'b11100_011101_00101;
        tomato_rice[22][19] = 16'b11011_011001_00100;
        tomato_rice[22][20] = 16'b11010_010010_00010;
        tomato_rice[22][21] = 16'b11011_010101_00010;
        tomato_rice[22][22] = 16'b11100_100000_00111;
        tomato_rice[22][23] = 16'b11110_110000_11110;
        tomato_rice[22][24] = 16'b11110_110000_11110;
        tomato_rice[22][25] = 16'b11110_110000_11110;
        tomato_rice[22][26] = 16'b11110_110000_11110;
        tomato_rice[22][27] = 16'b11110_110000_11110;
        tomato_rice[22][28] = 16'b11110_110000_11110;
        tomato_rice[22][29] = 16'b11110_110000_11110;
        tomato_rice[22][30] = 16'b11110_110000_11110;
        tomato_rice[22][31] = 16'b11110_110000_11110;
        tomato_rice[23][0] = 16'b11110_110000_11110;
        tomato_rice[23][1] = 16'b11110_110000_11110;
        tomato_rice[23][2] = 16'b11110_110000_11110;
        tomato_rice[23][3] = 16'b11110_110000_11110;
        tomato_rice[23][4] = 16'b11110_110000_11110;
        tomato_rice[23][5] = 16'b11110_110000_11110;
        tomato_rice[23][6] = 16'b11110_110000_11110;
        tomato_rice[23][7] = 16'b11110_110000_11110;
        tomato_rice[23][8] = 16'b11110_110000_11110;
        tomato_rice[23][9] = 16'b11110_110000_11110;
        tomato_rice[23][10] = 16'b11110_110000_11110;
        tomato_rice[23][11] = 16'b11100_100001_01000;
        tomato_rice[23][12] = 16'b11100_011010_00101;
        tomato_rice[23][13] = 16'b11011_010110_00011;
        tomato_rice[23][14] = 16'b11100_011001_00100;
        tomato_rice[23][15] = 16'b11011_010111_00011;
        tomato_rice[23][16] = 16'b11100_011001_00100;
        tomato_rice[23][17] = 16'b11100_011000_00100;
        tomato_rice[23][18] = 16'b11100_011000_00100;
        tomato_rice[23][19] = 16'b11011_010110_00011;
        tomato_rice[23][20] = 16'b11011_010110_00011;
        tomato_rice[23][21] = 16'b11110_110000_11110;
        tomato_rice[23][22] = 16'b11110_110000_11110;
        tomato_rice[23][23] = 16'b11110_110000_11110;
        tomato_rice[23][24] = 16'b11110_110000_11110;
        tomato_rice[23][25] = 16'b11110_110000_11110;
        tomato_rice[23][26] = 16'b11110_110000_11110;
        tomato_rice[23][27] = 16'b11110_110000_11110;
        tomato_rice[23][28] = 16'b11110_110000_11110;
        tomato_rice[23][29] = 16'b11110_110000_11110;
        tomato_rice[23][30] = 16'b11110_110000_11110;
        tomato_rice[23][31] = 16'b11110_110000_11110;
        tomato_rice[24][0] = 16'b11110_110000_11110;
        tomato_rice[24][1] = 16'b11110_110000_11110;
        tomato_rice[24][2] = 16'b11110_110000_11110;
        tomato_rice[24][3] = 16'b11110_110000_11110;
        tomato_rice[24][4] = 16'b11110_110000_11110;
        tomato_rice[24][5] = 16'b11110_110000_11110;
        tomato_rice[24][6] = 16'b11110_110000_11110;
        tomato_rice[24][7] = 16'b11110_110000_11110;
        tomato_rice[24][8] = 16'b11110_110000_11110;
        tomato_rice[24][9] = 16'b11110_110000_11110;
        tomato_rice[24][10] = 16'b11110_110000_11110;
        tomato_rice[24][11] = 16'b11110_110000_11110;
        tomato_rice[24][12] = 16'b11110_110000_11110;
        tomato_rice[24][13] = 16'b11100_011011_00101;
        tomato_rice[24][14] = 16'b11011_010101_00010;
        tomato_rice[24][15] = 16'b11100_011010_00100;
        tomato_rice[24][16] = 16'b11011_010101_00010;
        tomato_rice[24][17] = 16'b11100_011010_00100;
        tomato_rice[24][18] = 16'b11011_010101_00010;
        tomato_rice[24][19] = 16'b11110_110000_11110;
        tomato_rice[24][20] = 16'b11110_110000_11110;
        tomato_rice[24][21] = 16'b11110_110000_11110;
        tomato_rice[24][22] = 16'b11110_110000_11110;
        tomato_rice[24][23] = 16'b11110_110000_11110;
        tomato_rice[24][24] = 16'b11110_110000_11110;
        tomato_rice[24][25] = 16'b11110_110000_11110;
        tomato_rice[24][26] = 16'b11110_110000_11110;
        tomato_rice[24][27] = 16'b11110_110000_11110;
        tomato_rice[24][28] = 16'b11110_110000_11110;
        tomato_rice[24][29] = 16'b11110_110000_11110;
        tomato_rice[24][30] = 16'b11110_110000_11110;
        tomato_rice[24][31] = 16'b11110_110000_11110;
        tomato_rice[25][0] = 16'b11110_110000_11110;
        tomato_rice[25][1] = 16'b11110_110000_11110;
        tomato_rice[25][2] = 16'b11110_110000_11110;
        tomato_rice[25][3] = 16'b11110_110000_11110;
        tomato_rice[25][4] = 16'b11110_110000_11110;
        tomato_rice[25][5] = 16'b11110_110000_11110;
        tomato_rice[25][6] = 16'b11110_110000_11110;
        tomato_rice[25][7] = 16'b11110_110000_11110;
        tomato_rice[25][8] = 16'b11110_110000_11110;
        tomato_rice[25][9] = 16'b11110_110000_11110;
        tomato_rice[25][10] = 16'b11110_110000_11110;
        tomato_rice[25][11] = 16'b11110_110000_11110;
        tomato_rice[25][12] = 16'b11110_110000_11110;
        tomato_rice[25][13] = 16'b11110_110000_11110;
        tomato_rice[25][14] = 16'b11110_110000_11110;
        tomato_rice[25][15] = 16'b11110_110000_11110;
        tomato_rice[25][16] = 16'b11110_110000_11110;
        tomato_rice[25][17] = 16'b11110_110000_11110;
        tomato_rice[25][18] = 16'b11110_110000_11110;
        tomato_rice[25][19] = 16'b11110_110000_11110;
        tomato_rice[25][20] = 16'b11110_110000_11110;
        tomato_rice[25][21] = 16'b11110_110000_11110;
        tomato_rice[25][22] = 16'b11110_110000_11110;
        tomato_rice[25][23] = 16'b11110_110000_11110;
        tomato_rice[25][24] = 16'b11110_110000_11110;
        tomato_rice[25][25] = 16'b11110_110000_11110;
        tomato_rice[25][26] = 16'b11110_110000_11110;
        tomato_rice[25][27] = 16'b11110_110000_11110;
        tomato_rice[25][28] = 16'b11110_110000_11110;
        tomato_rice[25][29] = 16'b11110_110000_11110;
        tomato_rice[25][30] = 16'b11110_110000_11110;
        tomato_rice[25][31] = 16'b11110_110000_11110;
        tomato_rice[26][0] = 16'b11110_110000_11110;
        tomato_rice[26][1] = 16'b11110_110000_11110;
        tomato_rice[26][2] = 16'b11110_110000_11110;
        tomato_rice[26][3] = 16'b11110_110000_11110;
        tomato_rice[26][4] = 16'b11110_110000_11110;
        tomato_rice[26][5] = 16'b11110_110000_11110;
        tomato_rice[26][6] = 16'b11110_110000_11110;
        tomato_rice[26][7] = 16'b11110_110000_11110;
        tomato_rice[26][8] = 16'b11110_110000_11110;
        tomato_rice[26][9] = 16'b11110_110000_11110;
        tomato_rice[26][10] = 16'b11110_110000_11110;
        tomato_rice[26][11] = 16'b11110_110000_11110;
        tomato_rice[26][12] = 16'b11110_110000_11110;
        tomato_rice[26][13] = 16'b11110_110000_11110;
        tomato_rice[26][14] = 16'b11110_110000_11110;
        tomato_rice[26][15] = 16'b11110_110000_11110;
        tomato_rice[26][16] = 16'b11110_110000_11110;
        tomato_rice[26][17] = 16'b11110_110000_11110;
        tomato_rice[26][18] = 16'b11110_110000_11110;
        tomato_rice[26][19] = 16'b11110_110000_11110;
        tomato_rice[26][20] = 16'b11110_110000_11110;
        tomato_rice[26][21] = 16'b11110_110000_11110;
        tomato_rice[26][22] = 16'b11110_110000_11110;
        tomato_rice[26][23] = 16'b11110_110000_11110;
        tomato_rice[26][24] = 16'b11110_110000_11110;
        tomato_rice[26][25] = 16'b11110_110000_11110;
        tomato_rice[26][26] = 16'b11110_110000_11110;
        tomato_rice[26][27] = 16'b11110_110000_11110;
        tomato_rice[26][28] = 16'b11110_110000_11110;
        tomato_rice[26][29] = 16'b11110_110000_11110;
        tomato_rice[26][30] = 16'b11110_110000_11110;
        tomato_rice[26][31] = 16'b11110_110000_11110;
        tomato_rice[27][0] = 16'b11110_110000_11110;
        tomato_rice[27][1] = 16'b11110_110000_11110;
        tomato_rice[27][2] = 16'b11110_110000_11110;
        tomato_rice[27][3] = 16'b11110_110000_11110;
        tomato_rice[27][4] = 16'b11110_110000_11110;
        tomato_rice[27][5] = 16'b11110_110000_11110;
        tomato_rice[27][6] = 16'b11110_110000_11110;
        tomato_rice[27][7] = 16'b11110_110000_11110;
        tomato_rice[27][8] = 16'b11110_110000_11110;
        tomato_rice[27][9] = 16'b11110_110000_11110;
        tomato_rice[27][10] = 16'b11110_110000_11110;
        tomato_rice[27][11] = 16'b11110_110000_11110;
        tomato_rice[27][12] = 16'b11110_110000_11110;
        tomato_rice[27][13] = 16'b11110_110000_11110;
        tomato_rice[27][14] = 16'b11110_110000_11110;
        tomato_rice[27][15] = 16'b11110_110000_11110;
        tomato_rice[27][16] = 16'b11110_110000_11110;
        tomato_rice[27][17] = 16'b11110_110000_11110;
        tomato_rice[27][18] = 16'b11110_110000_11110;
        tomato_rice[27][19] = 16'b11110_110000_11110;
        tomato_rice[27][20] = 16'b11110_110000_11110;
        tomato_rice[27][21] = 16'b11110_110000_11110;
        tomato_rice[27][22] = 16'b11110_110000_11110;
        tomato_rice[27][23] = 16'b11110_110000_11110;
        tomato_rice[27][24] = 16'b11110_110000_11110;
        tomato_rice[27][25] = 16'b11110_110000_11110;
        tomato_rice[27][26] = 16'b11110_110000_11110;
        tomato_rice[27][27] = 16'b11110_110000_11110;
        tomato_rice[27][28] = 16'b11110_110000_11110;
        tomato_rice[27][29] = 16'b11110_110000_11110;
        tomato_rice[27][30] = 16'b11110_110000_11110;
        tomato_rice[27][31] = 16'b11110_110000_11110;
        tomato_rice[28][0] = 16'b11110_110000_11110;
        tomato_rice[28][1] = 16'b11110_110000_11110;
        tomato_rice[28][2] = 16'b11110_110000_11110;
        tomato_rice[28][3] = 16'b11110_110000_11110;
        tomato_rice[28][4] = 16'b11110_110000_11110;
        tomato_rice[28][5] = 16'b11110_110000_11110;
        tomato_rice[28][6] = 16'b11110_110000_11110;
        tomato_rice[28][7] = 16'b11110_110000_11110;
        tomato_rice[28][8] = 16'b11110_110000_11110;
        tomato_rice[28][9] = 16'b11110_110000_11110;
        tomato_rice[28][10] = 16'b11110_110000_11110;
        tomato_rice[28][11] = 16'b11110_110000_11110;
        tomato_rice[28][12] = 16'b11110_110000_11110;
        tomato_rice[28][13] = 16'b11110_110000_11110;
        tomato_rice[28][14] = 16'b11110_110000_11110;
        tomato_rice[28][15] = 16'b11110_110000_11110;
        tomato_rice[28][16] = 16'b11110_110000_11110;
        tomato_rice[28][17] = 16'b11110_110000_11110;
        tomato_rice[28][18] = 16'b11110_110000_11110;
        tomato_rice[28][19] = 16'b11110_110000_11110;
        tomato_rice[28][20] = 16'b11110_110000_11110;
        tomato_rice[28][21] = 16'b11110_110000_11110;
        tomato_rice[28][22] = 16'b11110_110000_11110;
        tomato_rice[28][23] = 16'b11110_110000_11110;
        tomato_rice[28][24] = 16'b11110_110000_11110;
        tomato_rice[28][25] = 16'b11110_110000_11110;
        tomato_rice[28][26] = 16'b11110_110000_11110;
        tomato_rice[28][27] = 16'b11110_110000_11110;
        tomato_rice[28][28] = 16'b11110_110000_11110;
        tomato_rice[28][29] = 16'b11110_110000_11110;
        tomato_rice[28][30] = 16'b11110_110000_11110;
        tomato_rice[28][31] = 16'b11110_110000_11110;
        tomato_rice[29][0] = 16'b11110_110000_11110;
        tomato_rice[29][1] = 16'b11110_110000_11110;
        tomato_rice[29][2] = 16'b11110_110000_11110;
        tomato_rice[29][3] = 16'b11110_110000_11110;
        tomato_rice[29][4] = 16'b11110_110000_11110;
        tomato_rice[29][5] = 16'b11110_110000_11110;
        tomato_rice[29][6] = 16'b11110_110000_11110;
        tomato_rice[29][7] = 16'b11110_110000_11110;
        tomato_rice[29][8] = 16'b11110_110000_11110;
        tomato_rice[29][9] = 16'b11110_110000_11110;
        tomato_rice[29][10] = 16'b11110_110000_11110;
        tomato_rice[29][11] = 16'b11110_110000_11110;
        tomato_rice[29][12] = 16'b11110_110000_11110;
        tomato_rice[29][13] = 16'b11110_110000_11110;
        tomato_rice[29][14] = 16'b11110_110000_11110;
        tomato_rice[29][15] = 16'b11110_110000_11110;
        tomato_rice[29][16] = 16'b11110_110000_11110;
        tomato_rice[29][17] = 16'b11110_110000_11110;
        tomato_rice[29][18] = 16'b11110_110000_11110;
        tomato_rice[29][19] = 16'b11110_110000_11110;
        tomato_rice[29][20] = 16'b11110_110000_11110;
        tomato_rice[29][21] = 16'b11110_110000_11110;
        tomato_rice[29][22] = 16'b11110_110000_11110;
        tomato_rice[29][23] = 16'b11110_110000_11110;
        tomato_rice[29][24] = 16'b11110_110000_11110;
        tomato_rice[29][25] = 16'b11110_110000_11110;
        tomato_rice[29][26] = 16'b11110_110000_11110;
        tomato_rice[29][27] = 16'b11110_110000_11110;
        tomato_rice[29][28] = 16'b11110_110000_11110;
        tomato_rice[29][29] = 16'b11110_110000_11110;
        tomato_rice[29][30] = 16'b11110_110000_11110;
        tomato_rice[29][31] = 16'b11110_110000_11110;
        tomato_rice[30][0] = 16'b11110_110000_11110;
        tomato_rice[30][1] = 16'b11110_110000_11110;
        tomato_rice[30][2] = 16'b11110_110000_11110;
        tomato_rice[30][3] = 16'b11110_110000_11110;
        tomato_rice[30][4] = 16'b11110_110000_11110;
        tomato_rice[30][5] = 16'b11110_110000_11110;
        tomato_rice[30][6] = 16'b11110_110000_11110;
        tomato_rice[30][7] = 16'b11110_110000_11110;
        tomato_rice[30][8] = 16'b11110_110000_11110;
        tomato_rice[30][9] = 16'b11110_110000_11110;
        tomato_rice[30][10] = 16'b11110_110000_11110;
        tomato_rice[30][11] = 16'b11110_110000_11110;
        tomato_rice[30][12] = 16'b11110_110000_11110;
        tomato_rice[30][13] = 16'b11110_110000_11110;
        tomato_rice[30][14] = 16'b11110_110000_11110;
        tomato_rice[30][15] = 16'b11110_110000_11110;
        tomato_rice[30][16] = 16'b11110_110000_11110;
        tomato_rice[30][17] = 16'b11110_110000_11110;
        tomato_rice[30][18] = 16'b11110_110000_11110;
        tomato_rice[30][19] = 16'b11110_110000_11110;
        tomato_rice[30][20] = 16'b11110_110000_11110;
        tomato_rice[30][21] = 16'b11110_110000_11110;
        tomato_rice[30][22] = 16'b11110_110000_11110;
        tomato_rice[30][23] = 16'b11110_110000_11110;
        tomato_rice[30][24] = 16'b11110_110000_11110;
        tomato_rice[30][25] = 16'b11110_110000_11110;
        tomato_rice[30][26] = 16'b11110_110000_11110;
        tomato_rice[30][27] = 16'b11110_110000_11110;
        tomato_rice[30][28] = 16'b11110_110000_11110;
        tomato_rice[30][29] = 16'b11110_110000_11110;
        tomato_rice[30][30] = 16'b11110_110000_11110;
        tomato_rice[30][31] = 16'b11110_110000_11110;
        tomato_rice[31][0] = 16'b11110_110000_11110;
        tomato_rice[31][1] = 16'b11110_110000_11110;
        tomato_rice[31][2] = 16'b11110_110000_11110;
        tomato_rice[31][3] = 16'b11110_110000_11110;
        tomato_rice[31][4] = 16'b11110_110000_11110;
        tomato_rice[31][5] = 16'b11110_110000_11110;
        tomato_rice[31][6] = 16'b11110_110000_11110;
        tomato_rice[31][7] = 16'b11110_110000_11110;
        tomato_rice[31][8] = 16'b11110_110000_11110;
        tomato_rice[31][9] = 16'b11110_110000_11110;
        tomato_rice[31][10] = 16'b11110_110000_11110;
        tomato_rice[31][11] = 16'b11110_110000_11110;
        tomato_rice[31][12] = 16'b11110_110000_11110;
        tomato_rice[31][13] = 16'b11110_110000_11110;
        tomato_rice[31][14] = 16'b11110_110000_11110;
        tomato_rice[31][15] = 16'b11110_110000_11110;
        tomato_rice[31][16] = 16'b11110_110000_11110;
        tomato_rice[31][17] = 16'b11110_110000_11110;
        tomato_rice[31][18] = 16'b11110_110000_11110;
        tomato_rice[31][19] = 16'b11110_110000_11110;
        tomato_rice[31][20] = 16'b11110_110000_11110;
        tomato_rice[31][21] = 16'b11110_110000_11110;
        tomato_rice[31][22] = 16'b11110_110000_11110;
        tomato_rice[31][23] = 16'b11110_110000_11110;
        tomato_rice[31][24] = 16'b11110_110000_11110;
        tomato_rice[31][25] = 16'b11110_110000_11110;
        tomato_rice[31][26] = 16'b11110_110000_11110;
        tomato_rice[31][27] = 16'b11110_110000_11110;
        tomato_rice[31][28] = 16'b11110_110000_11110;
        tomato_rice[31][29] = 16'b11110_110000_11110;
        tomato_rice[31][30] = 16'b11110_110000_11110;
        tomato_rice[31][31] = 16'b11110_110000_11110;
        
        chicken_rice_dim[0][0] = 16'b01011_011011_01111;
        chicken_rice_dim[0][1] = 16'b01011_011011_01111;
        chicken_rice_dim[0][2] = 16'b01011_011011_01111;
        chicken_rice_dim[0][3] = 16'b01011_011011_01111;
        chicken_rice_dim[0][4] = 16'b01011_011011_01111;
        chicken_rice_dim[0][5] = 16'b01011_011011_01111;
        chicken_rice_dim[0][6] = 16'b01011_011011_01111;
        chicken_rice_dim[0][7] = 16'b01011_011011_01111;
        chicken_rice_dim[0][8] = 16'b01011_011011_01111;
        chicken_rice_dim[0][9] = 16'b01011_011011_01111;
        chicken_rice_dim[0][10] = 16'b01011_011011_01111;
        chicken_rice_dim[0][11] = 16'b01011_011011_01111;
        chicken_rice_dim[0][12] = 16'b01011_011011_01111;
        chicken_rice_dim[0][13] = 16'b01011_011011_01111;
        chicken_rice_dim[0][14] = 16'b01011_011011_01111;
        chicken_rice_dim[0][15] = 16'b01011_011011_01111;
        chicken_rice_dim[0][16] = 16'b01011_011011_01111;
        chicken_rice_dim[0][17] = 16'b01011_011011_01111;
        chicken_rice_dim[0][18] = 16'b01011_011011_01111;
        chicken_rice_dim[0][19] = 16'b01011_011011_01111;
        chicken_rice_dim[0][20] = 16'b01011_011011_01111;
        chicken_rice_dim[0][21] = 16'b01011_011011_01111;
        chicken_rice_dim[0][22] = 16'b01011_011011_01111;
        chicken_rice_dim[0][23] = 16'b01011_011011_01111;
        chicken_rice_dim[0][24] = 16'b01011_011011_01111;
        chicken_rice_dim[0][25] = 16'b01011_011011_01111;
        chicken_rice_dim[0][26] = 16'b01011_011011_01111;
        chicken_rice_dim[0][27] = 16'b01011_011011_01111;
        chicken_rice_dim[0][28] = 16'b01011_011011_01111;
        chicken_rice_dim[0][29] = 16'b01011_011011_01111;
        chicken_rice_dim[0][30] = 16'b01011_011011_01111;
        chicken_rice_dim[0][31] = 16'b01011_011011_01111;
        chicken_rice_dim[1][0] = 16'b01011_011011_01111;
        chicken_rice_dim[1][1] = 16'b01011_011011_01111;
        chicken_rice_dim[1][2] = 16'b01011_011011_01111;
        chicken_rice_dim[1][3] = 16'b01011_011011_01111;
        chicken_rice_dim[1][4] = 16'b01011_011011_01111;
        chicken_rice_dim[1][5] = 16'b01011_011011_01111;
        chicken_rice_dim[1][6] = 16'b01011_011011_01111;
        chicken_rice_dim[1][7] = 16'b01011_011011_01111;
        chicken_rice_dim[1][8] = 16'b01011_011011_01111;
        chicken_rice_dim[1][9] = 16'b01011_011011_01111;
        chicken_rice_dim[1][10] = 16'b01011_011011_01111;
        chicken_rice_dim[1][11] = 16'b01011_011011_01111;
        chicken_rice_dim[1][12] = 16'b01011_011011_01111;
        chicken_rice_dim[1][13] = 16'b01011_011011_01111;
        chicken_rice_dim[1][14] = 16'b01011_011011_01111;
        chicken_rice_dim[1][15] = 16'b01011_011011_01111;
        chicken_rice_dim[1][16] = 16'b01011_011011_01111;
        chicken_rice_dim[1][17] = 16'b01011_011011_01111;
        chicken_rice_dim[1][18] = 16'b01011_011011_01111;
        chicken_rice_dim[1][19] = 16'b01011_011011_01111;
        chicken_rice_dim[1][20] = 16'b01011_011011_01111;
        chicken_rice_dim[1][21] = 16'b01011_011011_01111;
        chicken_rice_dim[1][22] = 16'b01011_011011_01111;
        chicken_rice_dim[1][23] = 16'b01011_011011_01111;
        chicken_rice_dim[1][24] = 16'b01011_011011_01111;
        chicken_rice_dim[1][25] = 16'b01011_011011_01111;
        chicken_rice_dim[1][26] = 16'b01011_011011_01111;
        chicken_rice_dim[1][27] = 16'b01011_011011_01111;
        chicken_rice_dim[1][28] = 16'b01011_011011_01111;
        chicken_rice_dim[1][29] = 16'b01011_011011_01111;
        chicken_rice_dim[1][30] = 16'b01011_011011_01111;
        chicken_rice_dim[1][31] = 16'b01011_011011_01111;
        chicken_rice_dim[2][0] = 16'b01011_011011_01111;
        chicken_rice_dim[2][1] = 16'b01011_011011_01111;
        chicken_rice_dim[2][2] = 16'b01011_011011_01111;
        chicken_rice_dim[2][3] = 16'b01011_011011_01111;
        chicken_rice_dim[2][4] = 16'b01011_011011_01111;
        chicken_rice_dim[2][5] = 16'b01011_011011_01111;
        chicken_rice_dim[2][6] = 16'b01011_011011_01111;
        chicken_rice_dim[2][7] = 16'b01011_011011_01111;
        chicken_rice_dim[2][8] = 16'b01011_011011_01111;
        chicken_rice_dim[2][9] = 16'b01011_011011_01111;
        chicken_rice_dim[2][10] = 16'b01011_011011_01111;
        chicken_rice_dim[2][11] = 16'b01011_011011_01111;
        chicken_rice_dim[2][12] = 16'b01011_011011_01111;
        chicken_rice_dim[2][13] = 16'b01011_011011_01111;
        chicken_rice_dim[2][14] = 16'b01011_011011_01111;
        chicken_rice_dim[2][15] = 16'b01011_011011_01111;
        chicken_rice_dim[2][16] = 16'b01011_011011_01111;
        chicken_rice_dim[2][17] = 16'b01011_011011_01111;
        chicken_rice_dim[2][18] = 16'b01011_011011_01111;
        chicken_rice_dim[2][19] = 16'b01011_011011_01111;
        chicken_rice_dim[2][20] = 16'b01011_011011_01111;
        chicken_rice_dim[2][21] = 16'b01011_011011_01111;
        chicken_rice_dim[2][22] = 16'b01011_011011_01111;
        chicken_rice_dim[2][23] = 16'b01011_011011_01111;
        chicken_rice_dim[2][24] = 16'b01011_011011_01111;
        chicken_rice_dim[2][25] = 16'b01011_011011_01111;
        chicken_rice_dim[2][26] = 16'b01011_011011_01111;
        chicken_rice_dim[2][27] = 16'b01011_011011_01111;
        chicken_rice_dim[2][28] = 16'b01011_011011_01111;
        chicken_rice_dim[2][29] = 16'b01011_011011_01111;
        chicken_rice_dim[2][30] = 16'b01011_011011_01111;
        chicken_rice_dim[2][31] = 16'b01011_011011_01111;
        chicken_rice_dim[3][0] = 16'b01011_011011_01111;
        chicken_rice_dim[3][1] = 16'b01011_011011_01111;
        chicken_rice_dim[3][2] = 16'b01011_011011_01111;
        chicken_rice_dim[3][3] = 16'b01011_011011_01111;
        chicken_rice_dim[3][4] = 16'b01011_011011_01111;
        chicken_rice_dim[3][5] = 16'b01011_011011_01111;
        chicken_rice_dim[3][6] = 16'b01011_011011_01111;
        chicken_rice_dim[3][7] = 16'b01011_011011_01111;
        chicken_rice_dim[3][8] = 16'b01011_011011_01111;
        chicken_rice_dim[3][9] = 16'b01011_011011_01111;
        chicken_rice_dim[3][10] = 16'b01011_011011_01111;
        chicken_rice_dim[3][11] = 16'b01011_011011_01111;
        chicken_rice_dim[3][12] = 16'b01011_011011_01111;
        chicken_rice_dim[3][13] = 16'b01011_011011_01111;
        chicken_rice_dim[3][14] = 16'b01011_011011_01111;
        chicken_rice_dim[3][15] = 16'b01011_011011_01111;
        chicken_rice_dim[3][16] = 16'b01011_011011_01111;
        chicken_rice_dim[3][17] = 16'b01011_011011_01111;
        chicken_rice_dim[3][18] = 16'b01011_011011_01111;
        chicken_rice_dim[3][19] = 16'b01011_011011_01111;
        chicken_rice_dim[3][20] = 16'b01011_011011_01111;
        chicken_rice_dim[3][21] = 16'b01011_011011_01111;
        chicken_rice_dim[3][22] = 16'b01011_011011_01111;
        chicken_rice_dim[3][23] = 16'b01011_011011_01111;
        chicken_rice_dim[3][24] = 16'b01011_011011_01111;
        chicken_rice_dim[3][25] = 16'b01011_011011_01111;
        chicken_rice_dim[3][26] = 16'b01011_011011_01111;
        chicken_rice_dim[3][27] = 16'b01011_011011_01111;
        chicken_rice_dim[3][28] = 16'b01011_011011_01111;
        chicken_rice_dim[3][29] = 16'b01011_011011_01111;
        chicken_rice_dim[3][30] = 16'b01011_011011_01111;
        chicken_rice_dim[3][31] = 16'b01011_011011_01111;
        chicken_rice_dim[4][0] = 16'b01011_011011_01111;
        chicken_rice_dim[4][1] = 16'b01011_011011_01111;
        chicken_rice_dim[4][2] = 16'b01011_011011_01111;
        chicken_rice_dim[4][3] = 16'b01011_011011_01111;
        chicken_rice_dim[4][4] = 16'b01011_011011_01111;
        chicken_rice_dim[4][5] = 16'b01011_011011_01111;
        chicken_rice_dim[4][6] = 16'b01011_011011_01111;
        chicken_rice_dim[4][7] = 16'b01011_011011_01111;
        chicken_rice_dim[4][8] = 16'b01011_011011_01111;
        chicken_rice_dim[4][9] = 16'b01011_011011_01111;
        chicken_rice_dim[4][10] = 16'b01011_011011_01111;
        chicken_rice_dim[4][11] = 16'b01011_011011_01111;
        chicken_rice_dim[4][12] = 16'b01011_011011_01111;
        chicken_rice_dim[4][13] = 16'b01011_011011_01111;
        chicken_rice_dim[4][14] = 16'b01011_011011_01111;
        chicken_rice_dim[4][15] = 16'b01011_011011_01111;
        chicken_rice_dim[4][16] = 16'b01011_011011_01111;
        chicken_rice_dim[4][17] = 16'b01011_011011_01111;
        chicken_rice_dim[4][18] = 16'b01011_011011_01111;
        chicken_rice_dim[4][19] = 16'b01011_011011_01111;
        chicken_rice_dim[4][20] = 16'b01011_011011_01111;
        chicken_rice_dim[4][21] = 16'b01011_011011_01111;
        chicken_rice_dim[4][22] = 16'b01011_011011_01111;
        chicken_rice_dim[4][23] = 16'b01011_011011_01111;
        chicken_rice_dim[4][24] = 16'b01011_011011_01111;
        chicken_rice_dim[4][25] = 16'b01011_011011_01111;
        chicken_rice_dim[4][26] = 16'b01011_011011_01111;
        chicken_rice_dim[4][27] = 16'b01011_011011_01111;
        chicken_rice_dim[4][28] = 16'b01011_011011_01111;
        chicken_rice_dim[4][29] = 16'b01011_011011_01111;
        chicken_rice_dim[4][30] = 16'b01011_011011_01111;
        chicken_rice_dim[4][31] = 16'b01011_011011_01111;
        chicken_rice_dim[5][0] = 16'b01011_011011_01111;
        chicken_rice_dim[5][1] = 16'b01011_011011_01111;
        chicken_rice_dim[5][2] = 16'b01011_011011_01111;
        chicken_rice_dim[5][3] = 16'b01011_011011_01111;
        chicken_rice_dim[5][4] = 16'b01011_011011_01111;
        chicken_rice_dim[5][5] = 16'b01011_011011_01111;
        chicken_rice_dim[5][6] = 16'b01011_011011_01111;
        chicken_rice_dim[5][7] = 16'b01011_011011_01111;
        chicken_rice_dim[5][8] = 16'b01011_011011_01111;
        chicken_rice_dim[5][9] = 16'b01011_011011_01111;
        chicken_rice_dim[5][10] = 16'b01011_011011_01111;
        chicken_rice_dim[5][11] = 16'b01011_011011_01111;
        chicken_rice_dim[5][12] = 16'b01100_010100_00110;
        chicken_rice_dim[5][13] = 16'b01101_010100_00110;
        chicken_rice_dim[5][14] = 16'b01101_010101_00110;
        chicken_rice_dim[5][15] = 16'b01101_010110_00111;
        chicken_rice_dim[5][16] = 16'b01101_010101_00111;
        chicken_rice_dim[5][17] = 16'b01110_011000_01000;
        chicken_rice_dim[5][18] = 16'b01101_010110_00111;
        chicken_rice_dim[5][19] = 16'b01011_011011_01111;
        chicken_rice_dim[5][20] = 16'b01011_011011_01111;
        chicken_rice_dim[5][21] = 16'b01011_011011_01111;
        chicken_rice_dim[5][22] = 16'b01011_011011_01111;
        chicken_rice_dim[5][23] = 16'b01011_011011_01111;
        chicken_rice_dim[5][24] = 16'b01011_011011_01111;
        chicken_rice_dim[5][25] = 16'b01011_011011_01111;
        chicken_rice_dim[5][26] = 16'b01011_011011_01111;
        chicken_rice_dim[5][27] = 16'b01011_011011_01111;
        chicken_rice_dim[5][28] = 16'b01011_011011_01111;
        chicken_rice_dim[5][29] = 16'b01011_011011_01111;
        chicken_rice_dim[5][30] = 16'b01011_011011_01111;
        chicken_rice_dim[5][31] = 16'b01011_011011_01111;
        chicken_rice_dim[6][0] = 16'b01011_011011_01111;
        chicken_rice_dim[6][1] = 16'b01011_011011_01111;
        chicken_rice_dim[6][2] = 16'b01011_011011_01111;
        chicken_rice_dim[6][3] = 16'b01011_011011_01111;
        chicken_rice_dim[6][4] = 16'b01011_011011_01111;
        chicken_rice_dim[6][5] = 16'b01011_011011_01111;
        chicken_rice_dim[6][6] = 16'b01011_011011_01111;
        chicken_rice_dim[6][7] = 16'b01011_011011_01111;
        chicken_rice_dim[6][8] = 16'b01011_011011_01111;
        chicken_rice_dim[6][9] = 16'b01100_010100_00110;
        chicken_rice_dim[6][10] = 16'b01110_010111_01000;
        chicken_rice_dim[6][11] = 16'b01101_010111_00111;
        chicken_rice_dim[6][12] = 16'b01101_010110_00111;
        chicken_rice_dim[6][13] = 16'b01101_010111_00111;
        chicken_rice_dim[6][14] = 16'b01110_010111_01000;
        chicken_rice_dim[6][15] = 16'b01110_011000_01000;
        chicken_rice_dim[6][16] = 16'b01110_010111_01000;
        chicken_rice_dim[6][17] = 16'b01110_011000_01000;
        chicken_rice_dim[6][18] = 16'b01110_011000_01000;
        chicken_rice_dim[6][19] = 16'b01110_011000_01000;
        chicken_rice_dim[6][20] = 16'b01110_011000_01000;
        chicken_rice_dim[6][21] = 16'b01110_011000_01000;
        chicken_rice_dim[6][22] = 16'b01101_010110_00111;
        chicken_rice_dim[6][23] = 16'b01011_011011_01111;
        chicken_rice_dim[6][24] = 16'b01011_011011_01111;
        chicken_rice_dim[6][25] = 16'b01011_011011_01111;
        chicken_rice_dim[6][26] = 16'b01011_011011_01111;
        chicken_rice_dim[6][27] = 16'b01011_011011_01111;
        chicken_rice_dim[6][28] = 16'b01011_011011_01111;
        chicken_rice_dim[6][29] = 16'b01011_011011_01111;
        chicken_rice_dim[6][30] = 16'b01011_011011_01111;
        chicken_rice_dim[6][31] = 16'b01011_011011_01111;
        chicken_rice_dim[7][0] = 16'b01011_011011_01111;
        chicken_rice_dim[7][1] = 16'b01011_011011_01111;
        chicken_rice_dim[7][2] = 16'b01011_011011_01111;
        chicken_rice_dim[7][3] = 16'b01011_011011_01111;
        chicken_rice_dim[7][4] = 16'b01011_011011_01111;
        chicken_rice_dim[7][5] = 16'b01011_011011_01111;
        chicken_rice_dim[7][6] = 16'b01011_011011_01111;
        chicken_rice_dim[7][7] = 16'b01100_010100_00110;
        chicken_rice_dim[7][8] = 16'b01110_010111_00111;
        chicken_rice_dim[7][9] = 16'b01101_010111_00111;
        chicken_rice_dim[7][10] = 16'b01101_010110_00111;
        chicken_rice_dim[7][11] = 16'b01101_010111_00111;
        chicken_rice_dim[7][12] = 16'b01101_010101_00111;
        chicken_rice_dim[7][13] = 16'b01101_010110_00111;
        chicken_rice_dim[7][14] = 16'b01101_010111_00111;
        chicken_rice_dim[7][15] = 16'b01101_010111_00111;
        chicken_rice_dim[7][16] = 16'b01101_010111_00111;
        chicken_rice_dim[7][17] = 16'b01101_010111_01000;
        chicken_rice_dim[7][18] = 16'b01110_011000_01000;
        chicken_rice_dim[7][19] = 16'b01110_011000_01000;
        chicken_rice_dim[7][20] = 16'b01110_011000_01000;
        chicken_rice_dim[7][21] = 16'b01110_011000_01000;
        chicken_rice_dim[7][22] = 16'b01110_011000_01000;
        chicken_rice_dim[7][23] = 16'b01110_011000_01000;
        chicken_rice_dim[7][24] = 16'b01011_011011_01111;
        chicken_rice_dim[7][25] = 16'b01011_011011_01111;
        chicken_rice_dim[7][26] = 16'b01011_011011_01111;
        chicken_rice_dim[7][27] = 16'b01011_011011_01111;
        chicken_rice_dim[7][28] = 16'b01011_011011_01111;
        chicken_rice_dim[7][29] = 16'b01011_011011_01111;
        chicken_rice_dim[7][30] = 16'b01011_011011_01111;
        chicken_rice_dim[7][31] = 16'b01011_011011_01111;
        chicken_rice_dim[8][0] = 16'b01011_011011_01111;
        chicken_rice_dim[8][1] = 16'b01011_011011_01111;
        chicken_rice_dim[8][2] = 16'b01011_011011_01111;
        chicken_rice_dim[8][3] = 16'b01011_011011_01111;
        chicken_rice_dim[8][4] = 16'b01011_011011_01111;
        chicken_rice_dim[8][5] = 16'b01011_011011_01111;
        chicken_rice_dim[8][6] = 16'b01100_010100_00110;
        chicken_rice_dim[8][7] = 16'b01101_010111_01000;
        chicken_rice_dim[8][8] = 16'b01101_010110_00111;
        chicken_rice_dim[8][9] = 16'b01011_001111_00011;
        chicken_rice_dim[8][10] = 16'b01011_001111_00011;
        chicken_rice_dim[8][11] = 16'b01100_010001_00100;
        chicken_rice_dim[8][12] = 16'b01100_010000_00011;
        chicken_rice_dim[8][13] = 16'b01100_010000_00011;
        chicken_rice_dim[8][14] = 16'b01100_010001_00011;
        chicken_rice_dim[8][15] = 16'b01011_001110_00010;
        chicken_rice_dim[8][16] = 16'b01100_010010_00100;
        chicken_rice_dim[8][17] = 16'b01100_010011_00101;
        chicken_rice_dim[8][18] = 16'b01100_010011_00101;
        chicken_rice_dim[8][19] = 16'b01100_010100_00110;
        chicken_rice_dim[8][20] = 16'b01101_010101_00110;
        chicken_rice_dim[8][21] = 16'b01101_010101_00110;
        chicken_rice_dim[8][22] = 16'b01101_010111_01000;
        chicken_rice_dim[8][23] = 16'b01110_011000_01000;
        chicken_rice_dim[8][24] = 16'b01110_011000_01000;
        chicken_rice_dim[8][25] = 16'b01101_010101_00110;
        chicken_rice_dim[8][26] = 16'b01011_011011_01111;
        chicken_rice_dim[8][27] = 16'b01011_011011_01111;
        chicken_rice_dim[8][28] = 16'b01011_011011_01111;
        chicken_rice_dim[8][29] = 16'b01011_011011_01111;
        chicken_rice_dim[8][30] = 16'b01011_011011_01111;
        chicken_rice_dim[8][31] = 16'b01011_011011_01111;
        chicken_rice_dim[9][0] = 16'b01011_011011_01111;
        chicken_rice_dim[9][1] = 16'b01011_011011_01111;
        chicken_rice_dim[9][2] = 16'b01011_011011_01111;
        chicken_rice_dim[9][3] = 16'b01011_011011_01111;
        chicken_rice_dim[9][4] = 16'b01100_010101_00111;
        chicken_rice_dim[9][5] = 16'b01110_011000_01000;
        chicken_rice_dim[9][6] = 16'b01110_011000_01000;
        chicken_rice_dim[9][7] = 16'b01100_010100_00110;
        chicken_rice_dim[9][8] = 16'b01011_001111_00010;
        chicken_rice_dim[9][9] = 16'b01011_001101_00001;
        chicken_rice_dim[9][10] = 16'b01100_001111_00001;
        chicken_rice_dim[9][11] = 16'b01101_010011_00011;
        chicken_rice_dim[9][12] = 16'b01110_010110_00110;
        chicken_rice_dim[9][13] = 16'b01110_011000_01000;
        chicken_rice_dim[9][14] = 16'b01101_010100_00101;
        chicken_rice_dim[9][15] = 16'b01100_010000_00010;
        chicken_rice_dim[9][16] = 16'b01011_001101_00010;
        chicken_rice_dim[9][17] = 16'b01011_010000_00011;
        chicken_rice_dim[9][18] = 16'b01100_010001_00100;
        chicken_rice_dim[9][19] = 16'b01100_010100_00110;
        chicken_rice_dim[9][20] = 16'b01100_010011_00101;
        chicken_rice_dim[9][21] = 16'b01100_010011_00101;
        chicken_rice_dim[9][22] = 16'b01100_010001_00100;
        chicken_rice_dim[9][23] = 16'b01100_010001_00100;
        chicken_rice_dim[9][24] = 16'b01110_010111_01000;
        chicken_rice_dim[9][25] = 16'b01101_010111_01000;
        chicken_rice_dim[9][26] = 16'b01110_010111_01000;
        chicken_rice_dim[9][27] = 16'b01100_010101_00110;
        chicken_rice_dim[9][28] = 16'b01011_011011_01111;
        chicken_rice_dim[9][29] = 16'b01011_011011_01111;
        chicken_rice_dim[9][30] = 16'b01011_011011_01111;
        chicken_rice_dim[9][31] = 16'b01011_011011_01111;
        chicken_rice_dim[10][0] = 16'b01011_011011_01111;
        chicken_rice_dim[10][1] = 16'b01011_011011_01111;
        chicken_rice_dim[10][2] = 16'b01011_011011_01111;
        chicken_rice_dim[10][3] = 16'b01101_010111_01000;
        chicken_rice_dim[10][4] = 16'b01110_011000_01000;
        chicken_rice_dim[10][5] = 16'b01110_011000_01000;
        chicken_rice_dim[10][6] = 16'b01101_010101_00110;
        chicken_rice_dim[10][7] = 16'b01100_010000_00011;
        chicken_rice_dim[10][8] = 16'b01011_001101_00001;
        chicken_rice_dim[10][9] = 16'b01101_010000_00001;
        chicken_rice_dim[10][10] = 16'b01101_010000_00001;
        chicken_rice_dim[10][11] = 16'b01101_010001_00010;
        chicken_rice_dim[10][12] = 16'b01101_010000_00010;
        chicken_rice_dim[10][13] = 16'b01101_010011_00100;
        chicken_rice_dim[10][14] = 16'b01110_010101_00101;
        chicken_rice_dim[10][15] = 16'b01101_010100_00101;
        chicken_rice_dim[10][16] = 16'b01100_001111_00010;
        chicken_rice_dim[10][17] = 16'b01100_010010_00100;
        chicken_rice_dim[10][18] = 16'b01101_010100_00101;
        chicken_rice_dim[10][19] = 16'b01110_011000_01000;
        chicken_rice_dim[10][20] = 16'b01101_010101_00110;
        chicken_rice_dim[10][21] = 16'b01101_010101_00110;
        chicken_rice_dim[10][22] = 16'b01101_010110_00111;
        chicken_rice_dim[10][23] = 16'b01101_010110_00111;
        chicken_rice_dim[10][24] = 16'b01100_010010_00100;
        chicken_rice_dim[10][25] = 16'b01101_010101_00110;
        chicken_rice_dim[10][26] = 16'b01110_010111_01000;
        chicken_rice_dim[10][27] = 16'b01110_011000_01000;
        chicken_rice_dim[10][28] = 16'b01101_010110_00111;
        chicken_rice_dim[10][29] = 16'b01011_011011_01111;
        chicken_rice_dim[10][30] = 16'b01011_011011_01111;
        chicken_rice_dim[10][31] = 16'b01011_011011_01111;
        chicken_rice_dim[11][0] = 16'b01011_011011_01111;
        chicken_rice_dim[11][1] = 16'b01011_011011_01111;
        chicken_rice_dim[11][2] = 16'b01011_011011_01111;
        chicken_rice_dim[11][3] = 16'b01110_011000_01000;
        chicken_rice_dim[11][4] = 16'b01110_011000_01000;
        chicken_rice_dim[11][5] = 16'b01110_011000_01000;
        chicken_rice_dim[11][6] = 16'b01100_010001_00100;
        chicken_rice_dim[11][7] = 16'b01011_001101_00001;
        chicken_rice_dim[11][8] = 16'b01100_001101_00000;
        chicken_rice_dim[11][9] = 16'b01110_010010_00010;
        chicken_rice_dim[11][10] = 16'b01110_010010_00010;
        chicken_rice_dim[11][11] = 16'b01110_010011_00010;
        chicken_rice_dim[11][12] = 16'b01110_010011_00011;
        chicken_rice_dim[11][13] = 16'b01110_010100_00100;
        chicken_rice_dim[11][14] = 16'b01100_010001_00011;
        chicken_rice_dim[11][15] = 16'b01101_010100_00101;
        chicken_rice_dim[11][16] = 16'b01101_010011_00100;
        chicken_rice_dim[11][17] = 16'b01100_010001_00100;
        chicken_rice_dim[11][18] = 16'b01101_010111_00111;
        chicken_rice_dim[11][19] = 16'b01110_011000_01000;
        chicken_rice_dim[11][20] = 16'b01110_011000_01000;
        chicken_rice_dim[11][21] = 16'b01101_010111_00111;
        chicken_rice_dim[11][22] = 16'b01110_011000_01000;
        chicken_rice_dim[11][23] = 16'b01110_011001_01000;
        chicken_rice_dim[11][24] = 16'b01101_010110_00111;
        chicken_rice_dim[11][25] = 16'b01011_010001_00100;
        chicken_rice_dim[11][26] = 16'b01101_010101_00111;
        chicken_rice_dim[11][27] = 16'b01101_010111_01000;
        chicken_rice_dim[11][28] = 16'b01110_011000_01000;
        chicken_rice_dim[11][29] = 16'b01011_011011_01111;
        chicken_rice_dim[11][30] = 16'b01011_011011_01111;
        chicken_rice_dim[11][31] = 16'b01011_011011_01111;
        chicken_rice_dim[12][0] = 16'b01011_011011_01111;
        chicken_rice_dim[12][1] = 16'b01011_011011_01111;
        chicken_rice_dim[12][2] = 16'b01101_010111_01000;
        chicken_rice_dim[12][3] = 16'b01110_011000_01000;
        chicken_rice_dim[12][4] = 16'b01110_011000_01000;
        chicken_rice_dim[12][5] = 16'b01101_010100_00110;
        chicken_rice_dim[12][6] = 16'b01100_001110_00010;
        chicken_rice_dim[12][7] = 16'b01101_001110_00000;
        chicken_rice_dim[12][8] = 16'b01100_001110_00000;
        chicken_rice_dim[12][9] = 16'b01100_001100_00000;
        chicken_rice_dim[12][10] = 16'b01110_010011_00010;
        chicken_rice_dim[12][11] = 16'b01110_010100_00100;
        chicken_rice_dim[12][12] = 16'b01110_010110_00101;
        chicken_rice_dim[12][13] = 16'b01110_010101_00100;
        chicken_rice_dim[12][14] = 16'b01101_010011_00011;
        chicken_rice_dim[12][15] = 16'b01101_010010_00011;
        chicken_rice_dim[12][16] = 16'b01101_010000_00010;
        chicken_rice_dim[12][17] = 16'b01011_001111_00011;
        chicken_rice_dim[12][18] = 16'b01101_010110_00110;
        chicken_rice_dim[12][19] = 16'b01110_011000_01000;
        chicken_rice_dim[12][20] = 16'b01110_011001_01001;
        chicken_rice_dim[12][21] = 16'b01101_010111_01000;
        chicken_rice_dim[12][22] = 16'b01101_010111_01000;
        chicken_rice_dim[12][23] = 16'b01110_011001_01001;
        chicken_rice_dim[12][24] = 16'b01110_011001_01000;
        chicken_rice_dim[12][25] = 16'b01101_010101_00110;
        chicken_rice_dim[12][26] = 16'b01100_010001_00100;
        chicken_rice_dim[12][27] = 16'b01101_010111_00111;
        chicken_rice_dim[12][28] = 16'b01110_011000_01000;
        chicken_rice_dim[12][29] = 16'b01110_011000_01000;
        chicken_rice_dim[12][30] = 16'b01011_011011_01111;
        chicken_rice_dim[12][31] = 16'b01011_011011_01111;
        chicken_rice_dim[13][0] = 16'b01011_011011_01111;
        chicken_rice_dim[13][1] = 16'b01011_011011_01111;
        chicken_rice_dim[13][2] = 16'b01110_011001_01001;
        chicken_rice_dim[13][3] = 16'b01110_011000_01000;
        chicken_rice_dim[13][4] = 16'b01110_011000_01000;
        chicken_rice_dim[13][5] = 16'b01100_010100_00101;
        chicken_rice_dim[13][6] = 16'b01011_001100_00000;
        chicken_rice_dim[13][7] = 16'b01101_010000_00001;
        chicken_rice_dim[13][8] = 16'b01101_010001_00001;
        chicken_rice_dim[13][9] = 16'b01011_001011_00000;
        chicken_rice_dim[13][10] = 16'b01011_001100_00000;
        chicken_rice_dim[13][11] = 16'b01101_010001_00001;
        chicken_rice_dim[13][12] = 16'b01101_010010_00010;
        chicken_rice_dim[13][13] = 16'b01110_010101_00101;
        chicken_rice_dim[13][14] = 16'b01101_010010_00010;
        chicken_rice_dim[13][15] = 16'b01101_010001_00010;
        chicken_rice_dim[13][16] = 16'b01101_001111_00001;
        chicken_rice_dim[13][17] = 16'b01100_001101_00000;
        chicken_rice_dim[13][18] = 16'b01110_010111_01000;
        chicken_rice_dim[13][19] = 16'b01110_011001_01001;
        chicken_rice_dim[13][20] = 16'b01110_011000_01000;
        chicken_rice_dim[13][21] = 16'b01101_010111_01000;
        chicken_rice_dim[13][22] = 16'b01110_011001_01001;
        chicken_rice_dim[13][23] = 16'b01110_011010_01001;
        chicken_rice_dim[13][24] = 16'b01110_011001_01000;
        chicken_rice_dim[13][25] = 16'b01110_011000_01000;
        chicken_rice_dim[13][26] = 16'b01100_010011_00101;
        chicken_rice_dim[13][27] = 16'b01101_010110_00111;
        chicken_rice_dim[13][28] = 16'b01110_011000_01000;
        chicken_rice_dim[13][29] = 16'b01110_011001_01000;
        chicken_rice_dim[13][30] = 16'b01011_011011_01111;
        chicken_rice_dim[13][31] = 16'b01011_011011_01111;
        chicken_rice_dim[14][0] = 16'b01011_011011_01111;
        chicken_rice_dim[14][1] = 16'b01011_011011_01111;
        chicken_rice_dim[14][2] = 16'b01110_011001_01001;
        chicken_rice_dim[14][3] = 16'b01110_011000_01000;
        chicken_rice_dim[14][4] = 16'b01101_010111_00111;
        chicken_rice_dim[14][5] = 16'b01011_001100_00001;
        chicken_rice_dim[14][6] = 16'b01010_001011_00000;
        chicken_rice_dim[14][7] = 16'b01011_001100_00000;
        chicken_rice_dim[14][8] = 16'b01101_010001_00001;
        chicken_rice_dim[14][9] = 16'b01110_010011_00010;
        chicken_rice_dim[14][10] = 16'b01110_010010_00010;
        chicken_rice_dim[14][11] = 16'b01100_001110_00000;
        chicken_rice_dim[14][12] = 16'b01100_001111_00000;
        chicken_rice_dim[14][13] = 16'b01101_010001_00010;
        chicken_rice_dim[14][14] = 16'b01110_010100_00011;
        chicken_rice_dim[14][15] = 16'b01110_010011_00011;
        chicken_rice_dim[14][16] = 16'b01110_010011_00011;
        chicken_rice_dim[14][17] = 16'b01101_010001_00010;
        chicken_rice_dim[14][18] = 16'b01101_010101_00111;
        chicken_rice_dim[14][19] = 16'b01110_011000_01000;
        chicken_rice_dim[14][20] = 16'b01110_011000_01000;
        chicken_rice_dim[14][21] = 16'b01110_011000_01000;
        chicken_rice_dim[14][22] = 16'b01110_011010_01001;
        chicken_rice_dim[14][23] = 16'b01110_011001_01001;
        chicken_rice_dim[14][24] = 16'b01110_011010_01001;
        chicken_rice_dim[14][25] = 16'b01110_011001_01001;
        chicken_rice_dim[14][26] = 16'b01101_010111_00111;
        chicken_rice_dim[14][27] = 16'b01100_010011_00101;
        chicken_rice_dim[14][28] = 16'b01110_011000_01000;
        chicken_rice_dim[14][29] = 16'b01110_011000_01000;
        chicken_rice_dim[14][30] = 16'b01011_011011_01111;
        chicken_rice_dim[14][31] = 16'b01011_011011_01111;
        chicken_rice_dim[15][0] = 16'b01011_011011_01111;
        chicken_rice_dim[15][1] = 16'b01011_011011_01111;
        chicken_rice_dim[15][2] = 16'b01110_011001_01001;
        chicken_rice_dim[15][3] = 16'b01110_011001_01000;
        chicken_rice_dim[15][4] = 16'b01101_010110_00111;
        chicken_rice_dim[15][5] = 16'b01011_001100_00000;
        chicken_rice_dim[15][6] = 16'b01101_001111_00000;
        chicken_rice_dim[15][7] = 16'b01011_001011_00000;
        chicken_rice_dim[15][8] = 16'b01100_001110_00001;
        chicken_rice_dim[15][9] = 16'b01110_010101_00011;
        chicken_rice_dim[15][10] = 16'b01110_010111_00101;
        chicken_rice_dim[15][11] = 16'b01110_010100_00100;
        chicken_rice_dim[15][12] = 16'b01110_010011_00011;
        chicken_rice_dim[15][13] = 16'b01101_010001_00010;
        chicken_rice_dim[15][14] = 16'b01101_010001_00010;
        chicken_rice_dim[15][15] = 16'b01100_001110_00001;
        chicken_rice_dim[15][16] = 16'b01100_001110_00001;
        chicken_rice_dim[15][17] = 16'b01101_010001_00010;
        chicken_rice_dim[15][18] = 16'b01101_010111_00111;
        chicken_rice_dim[15][19] = 16'b01110_011001_01001;
        chicken_rice_dim[15][20] = 16'b01110_011010_01010;
        chicken_rice_dim[15][21] = 16'b01110_011001_01001;
        chicken_rice_dim[15][22] = 16'b01110_011010_01001;
        chicken_rice_dim[15][23] = 16'b01110_011011_01010;
        chicken_rice_dim[15][24] = 16'b01110_011001_01001;
        chicken_rice_dim[15][25] = 16'b01110_011010_01001;
        chicken_rice_dim[15][26] = 16'b01110_011000_01000;
        chicken_rice_dim[15][27] = 16'b01100_010011_00101;
        chicken_rice_dim[15][28] = 16'b01110_011000_01000;
        chicken_rice_dim[15][29] = 16'b01110_011001_01000;
        chicken_rice_dim[15][30] = 16'b01011_011011_01111;
        chicken_rice_dim[15][31] = 16'b01011_011011_01111;
        chicken_rice_dim[16][0] = 16'b01011_011011_01111;
        chicken_rice_dim[16][1] = 16'b01011_011011_01111;
        chicken_rice_dim[16][2] = 16'b01110_011001_01001;
        chicken_rice_dim[16][3] = 16'b01110_011000_01000;
        chicken_rice_dim[16][4] = 16'b01101_010101_00110;
        chicken_rice_dim[16][5] = 16'b01011_001100_00001;
        chicken_rice_dim[16][6] = 16'b01101_010000_00001;
        chicken_rice_dim[16][7] = 16'b01101_010010_00010;
        chicken_rice_dim[16][8] = 16'b01101_001111_00000;
        chicken_rice_dim[16][9] = 16'b01101_010000_00000;
        chicken_rice_dim[16][10] = 16'b01110_010100_00011;
        chicken_rice_dim[16][11] = 16'b01110_011000_00111;
        chicken_rice_dim[16][12] = 16'b01110_011000_00111;
        chicken_rice_dim[16][13] = 16'b01110_010101_00100;
        chicken_rice_dim[16][14] = 16'b01101_010011_00011;
        chicken_rice_dim[16][15] = 16'b01100_001111_00000;
        chicken_rice_dim[16][16] = 16'b01100_001101_00000;
        chicken_rice_dim[16][17] = 16'b01110_010011_00011;
        chicken_rice_dim[16][18] = 16'b01110_011001_01001;
        chicken_rice_dim[16][19] = 16'b01110_011010_01001;
        chicken_rice_dim[16][20] = 16'b01110_011011_01010;
        chicken_rice_dim[16][21] = 16'b01110_011001_01001;
        chicken_rice_dim[16][22] = 16'b01110_011001_01001;
        chicken_rice_dim[16][23] = 16'b01111_011011_01010;
        chicken_rice_dim[16][24] = 16'b01110_011001_01001;
        chicken_rice_dim[16][25] = 16'b01110_011001_01001;
        chicken_rice_dim[16][26] = 16'b01110_011000_01000;
        chicken_rice_dim[16][27] = 16'b01100_010100_00101;
        chicken_rice_dim[16][28] = 16'b01110_011000_01000;
        chicken_rice_dim[16][29] = 16'b01110_011000_01000;
        chicken_rice_dim[16][30] = 16'b01011_011011_01111;
        chicken_rice_dim[16][31] = 16'b01011_011011_01111;
        chicken_rice_dim[17][0] = 16'b01011_011011_01111;
        chicken_rice_dim[17][1] = 16'b01011_011011_01111;
        chicken_rice_dim[17][2] = 16'b01110_011001_01001;
        chicken_rice_dim[17][3] = 16'b01110_011000_01000;
        chicken_rice_dim[17][4] = 16'b01101_010111_00111;
        chicken_rice_dim[17][5] = 16'b01011_001101_00000;
        chicken_rice_dim[17][6] = 16'b01101_010000_00001;
        chicken_rice_dim[17][7] = 16'b01110_010011_00011;
        chicken_rice_dim[17][8] = 16'b01110_010011_00011;
        chicken_rice_dim[17][9] = 16'b01101_010000_00000;
        chicken_rice_dim[17][10] = 16'b01101_001110_00000;
        chicken_rice_dim[17][11] = 16'b01101_010000_00001;
        chicken_rice_dim[17][12] = 16'b01101_010001_00010;
        chicken_rice_dim[17][13] = 16'b01101_010010_00011;
        chicken_rice_dim[17][14] = 16'b01101_010011_00011;
        chicken_rice_dim[17][15] = 16'b01100_001110_00000;
        chicken_rice_dim[17][16] = 16'b01011_001011_00000;
        chicken_rice_dim[17][17] = 16'b01110_010100_00011;
        chicken_rice_dim[17][18] = 16'b01110_011010_01001;
        chicken_rice_dim[17][19] = 16'b01111_011011_01010;
        chicken_rice_dim[17][20] = 16'b01110_011010_01001;
        chicken_rice_dim[17][21] = 16'b01111_011011_01010;
        chicken_rice_dim[17][22] = 16'b01110_011001_01001;
        chicken_rice_dim[17][23] = 16'b01110_011001_01001;
        chicken_rice_dim[17][24] = 16'b01110_011011_01010;
        chicken_rice_dim[17][25] = 16'b01110_011001_01001;
        chicken_rice_dim[17][26] = 16'b01101_010111_01000;
        chicken_rice_dim[17][27] = 16'b01100_010100_00110;
        chicken_rice_dim[17][28] = 16'b01101_011000_01000;
        chicken_rice_dim[17][29] = 16'b01110_011000_01000;
        chicken_rice_dim[17][30] = 16'b01011_011011_01111;
        chicken_rice_dim[17][31] = 16'b01011_011011_01111;
        chicken_rice_dim[18][0] = 16'b01011_011011_01111;
        chicken_rice_dim[18][1] = 16'b01011_011011_01111;
        chicken_rice_dim[18][2] = 16'b01110_011001_01001;
        chicken_rice_dim[18][3] = 16'b01110_011001_01000;
        chicken_rice_dim[18][4] = 16'b01110_011000_01000;
        chicken_rice_dim[18][5] = 16'b01101_010100_00101;
        chicken_rice_dim[18][6] = 16'b01100_001100_00000;
        chicken_rice_dim[18][7] = 16'b01100_001111_00001;
        chicken_rice_dim[18][8] = 16'b01110_010100_00011;
        chicken_rice_dim[18][9] = 16'b01110_010101_00101;
        chicken_rice_dim[18][10] = 16'b01110_010101_00100;
        chicken_rice_dim[18][11] = 16'b01101_010001_00010;
        chicken_rice_dim[18][12] = 16'b01100_001111_00001;
        chicken_rice_dim[18][13] = 16'b01101_010000_00001;
        chicken_rice_dim[18][14] = 16'b01011_001100_00000;
        chicken_rice_dim[18][15] = 16'b01011_001100_00000;
        chicken_rice_dim[18][16] = 16'b01100_001101_00000;
        chicken_rice_dim[18][17] = 16'b01110_011001_01001;
        chicken_rice_dim[18][18] = 16'b01110_011011_01010;
        chicken_rice_dim[18][19] = 16'b01110_011010_01001;
        chicken_rice_dim[18][20] = 16'b01110_011010_01001;
        chicken_rice_dim[18][21] = 16'b01110_011011_01010;
        chicken_rice_dim[18][22] = 16'b01110_011011_01010;
        chicken_rice_dim[18][23] = 16'b01110_011010_01001;
        chicken_rice_dim[18][24] = 16'b01110_011010_01001;
        chicken_rice_dim[18][25] = 16'b01110_011001_01001;
        chicken_rice_dim[18][26] = 16'b01101_010101_00110;
        chicken_rice_dim[18][27] = 16'b01101_010111_00111;
        chicken_rice_dim[18][28] = 16'b01110_011000_01000;
        chicken_rice_dim[18][29] = 16'b01110_011000_01000;
        chicken_rice_dim[18][30] = 16'b01011_011011_01111;
        chicken_rice_dim[18][31] = 16'b01011_011011_01111;
        chicken_rice_dim[19][0] = 16'b01011_011011_01111;
        chicken_rice_dim[19][1] = 16'b01011_011011_01111;
        chicken_rice_dim[19][2] = 16'b01011_011011_01111;
        chicken_rice_dim[19][3] = 16'b01110_011001_01001;
        chicken_rice_dim[19][4] = 16'b01110_011000_01000;
        chicken_rice_dim[19][5] = 16'b01110_011000_01000;
        chicken_rice_dim[19][6] = 16'b01101_010001_00010;
        chicken_rice_dim[19][7] = 16'b01100_001111_00001;
        chicken_rice_dim[19][8] = 16'b01100_010000_00001;
        chicken_rice_dim[19][9] = 16'b01110_010100_00100;
        chicken_rice_dim[19][10] = 16'b01110_010101_00101;
        chicken_rice_dim[19][11] = 16'b01110_010101_00100;
        chicken_rice_dim[19][12] = 16'b01110_010101_00100;
        chicken_rice_dim[19][13] = 16'b01101_010001_00010;
        chicken_rice_dim[19][14] = 16'b01101_010001_00010;
        chicken_rice_dim[19][15] = 16'b01100_001111_00001;
        chicken_rice_dim[19][16] = 16'b01101_010010_00010;
        chicken_rice_dim[19][17] = 16'b01110_011010_01010;
        chicken_rice_dim[19][18] = 16'b01110_011010_01001;
        chicken_rice_dim[19][19] = 16'b01110_011011_01010;
        chicken_rice_dim[19][20] = 16'b01110_011010_01001;
        chicken_rice_dim[19][21] = 16'b01110_011010_01001;
        chicken_rice_dim[19][22] = 16'b01110_011011_01010;
        chicken_rice_dim[19][23] = 16'b01110_011011_01010;
        chicken_rice_dim[19][24] = 16'b01110_011010_01010;
        chicken_rice_dim[19][25] = 16'b01110_011000_01000;
        chicken_rice_dim[19][26] = 16'b01101_010111_00111;
        chicken_rice_dim[19][27] = 16'b01101_010111_00111;
        chicken_rice_dim[19][28] = 16'b01110_011000_01000;
        chicken_rice_dim[19][29] = 16'b01011_011011_01111;
        chicken_rice_dim[19][30] = 16'b01011_011011_01111;
        chicken_rice_dim[19][31] = 16'b01011_011011_01111;
        chicken_rice_dim[20][0] = 16'b01011_011011_01111;
        chicken_rice_dim[20][1] = 16'b01011_011011_01111;
        chicken_rice_dim[20][2] = 16'b01011_011011_01111;
        chicken_rice_dim[20][3] = 16'b01110_011000_01000;
        chicken_rice_dim[20][4] = 16'b01110_011000_01000;
        chicken_rice_dim[20][5] = 16'b01110_011000_01000;
        chicken_rice_dim[20][6] = 16'b01110_010111_00111;
        chicken_rice_dim[20][7] = 16'b01101_010000_00001;
        chicken_rice_dim[20][8] = 16'b01101_010001_00001;
        chicken_rice_dim[20][9] = 16'b01101_010000_00001;
        chicken_rice_dim[20][10] = 16'b01101_010000_00001;
        chicken_rice_dim[20][11] = 16'b01101_010010_00010;
        chicken_rice_dim[20][12] = 16'b01101_010010_00010;
        chicken_rice_dim[20][13] = 16'b01101_010001_00010;
        chicken_rice_dim[20][14] = 16'b01100_001110_00000;
        chicken_rice_dim[20][15] = 16'b01100_001110_00000;
        chicken_rice_dim[20][16] = 16'b01110_011001_01001;
        chicken_rice_dim[20][17] = 16'b01111_011011_01010;
        chicken_rice_dim[20][18] = 16'b01110_011010_01001;
        chicken_rice_dim[20][19] = 16'b01111_011011_01010;
        chicken_rice_dim[20][20] = 16'b01111_011011_01010;
        chicken_rice_dim[20][21] = 16'b01110_011010_01001;
        chicken_rice_dim[20][22] = 16'b01110_011010_01010;
        chicken_rice_dim[20][23] = 16'b01110_011010_01001;
        chicken_rice_dim[20][24] = 16'b01110_011001_01001;
        chicken_rice_dim[20][25] = 16'b01001_010010_00101;
        chicken_rice_dim[20][26] = 16'b01101_010110_00111;
        chicken_rice_dim[20][27] = 16'b01101_010111_00111;
        chicken_rice_dim[20][28] = 16'b01101_011000_01000;
        chicken_rice_dim[20][29] = 16'b01011_011011_01111;
        chicken_rice_dim[20][30] = 16'b01011_011011_01111;
        chicken_rice_dim[20][31] = 16'b01011_011011_01111;
        chicken_rice_dim[21][0] = 16'b01011_011011_01111;
        chicken_rice_dim[21][1] = 16'b01011_011011_01111;
        chicken_rice_dim[21][2] = 16'b01011_011011_01111;
        chicken_rice_dim[21][3] = 16'b01011_011011_01111;
        chicken_rice_dim[21][4] = 16'b01101_010111_01000;
        chicken_rice_dim[21][5] = 16'b01110_011000_01000;
        chicken_rice_dim[21][6] = 16'b01110_011000_01000;
        chicken_rice_dim[21][7] = 16'b01101_010011_00101;
        chicken_rice_dim[21][8] = 16'b01101_010001_00010;
        chicken_rice_dim[21][9] = 16'b01110_010101_00100;
        chicken_rice_dim[21][10] = 16'b01110_010010_00010;
        chicken_rice_dim[21][11] = 16'b01101_010000_00001;
        chicken_rice_dim[21][12] = 16'b01100_001110_00001;
        chicken_rice_dim[21][13] = 16'b01011_001101_00000;
        chicken_rice_dim[21][14] = 16'b01100_001101_00000;
        chicken_rice_dim[21][15] = 16'b01101_010100_00110;
        chicken_rice_dim[21][16] = 16'b01111_011011_01010;
        chicken_rice_dim[21][17] = 16'b01111_011100_01011;
        chicken_rice_dim[21][18] = 16'b01111_011100_01011;
        chicken_rice_dim[21][19] = 16'b01111_011011_01010;
        chicken_rice_dim[21][20] = 16'b01110_011011_01010;
        chicken_rice_dim[21][21] = 16'b01111_011011_01010;
        chicken_rice_dim[21][22] = 16'b01111_011011_01010;
        chicken_rice_dim[21][23] = 16'b01110_011011_01010;
        chicken_rice_dim[21][24] = 16'b01001_010010_00101;
        chicken_rice_dim[21][25] = 16'b00110_001101_00010;
        chicken_rice_dim[21][26] = 16'b01101_010110_00111;
        chicken_rice_dim[21][27] = 16'b01101_010111_00111;
        chicken_rice_dim[21][28] = 16'b01011_011011_01111;
        chicken_rice_dim[21][29] = 16'b01011_011011_01111;
        chicken_rice_dim[21][30] = 16'b01011_011011_01111;
        chicken_rice_dim[21][31] = 16'b01011_011011_01111;
        chicken_rice_dim[22][0] = 16'b01011_011011_01111;
        chicken_rice_dim[22][1] = 16'b01011_011011_01111;
        chicken_rice_dim[22][2] = 16'b01011_011011_01111;
        chicken_rice_dim[22][3] = 16'b01011_011011_01111;
        chicken_rice_dim[22][4] = 16'b01011_011011_01111;
        chicken_rice_dim[22][5] = 16'b01101_010111_00111;
        chicken_rice_dim[22][6] = 16'b01101_010111_00111;
        chicken_rice_dim[22][7] = 16'b01101_010110_00111;
        chicken_rice_dim[22][8] = 16'b01101_010011_00100;
        chicken_rice_dim[22][9] = 16'b01110_010011_00011;
        chicken_rice_dim[22][10] = 16'b01110_010111_00110;
        chicken_rice_dim[22][11] = 16'b01110_010110_00101;
        chicken_rice_dim[22][12] = 16'b01101_010010_00100;
        chicken_rice_dim[22][13] = 16'b01101_010011_00100;
        chicken_rice_dim[22][14] = 16'b01100_001110_00000;
        chicken_rice_dim[22][15] = 16'b01100_010001_00100;
        chicken_rice_dim[22][16] = 16'b01111_011100_01011;
        chicken_rice_dim[22][17] = 16'b01111_011100_01011;
        chicken_rice_dim[22][18] = 16'b01111_011011_01010;
        chicken_rice_dim[22][19] = 16'b01111_011011_01010;
        chicken_rice_dim[22][20] = 16'b01110_011010_01010;
        chicken_rice_dim[22][21] = 16'b01110_011011_01010;
        chicken_rice_dim[22][22] = 16'b01111_011100_01011;
        chicken_rice_dim[22][23] = 16'b01110_011011_01010;
        chicken_rice_dim[22][24] = 16'b00111_001111_00011;
        chicken_rice_dim[22][25] = 16'b00110_001101_00010;
        chicken_rice_dim[22][26] = 16'b01100_010101_00111;
        chicken_rice_dim[22][27] = 16'b01011_011011_01111;
        chicken_rice_dim[22][28] = 16'b01011_011011_01111;
        chicken_rice_dim[22][29] = 16'b01011_011011_01111;
        chicken_rice_dim[22][30] = 16'b01011_011011_01111;
        chicken_rice_dim[22][31] = 16'b01011_011011_01111;
        chicken_rice_dim[23][0] = 16'b01011_011011_01111;
        chicken_rice_dim[23][1] = 16'b01011_011011_01111;
        chicken_rice_dim[23][2] = 16'b01011_011011_01111;
        chicken_rice_dim[23][3] = 16'b01011_011011_01111;
        chicken_rice_dim[23][4] = 16'b01011_011011_01111;
        chicken_rice_dim[23][5] = 16'b01011_011011_01111;
        chicken_rice_dim[23][6] = 16'b01011_011011_01111;
        chicken_rice_dim[23][7] = 16'b01011_011011_01111;
        chicken_rice_dim[23][8] = 16'b01110_011000_01000;
        chicken_rice_dim[23][9] = 16'b01110_011000_01000;
        chicken_rice_dim[23][10] = 16'b01110_011000_01000;
        chicken_rice_dim[23][11] = 16'b01110_011000_01000;
        chicken_rice_dim[23][12] = 16'b01110_011000_01000;
        chicken_rice_dim[23][13] = 16'b01110_011000_01000;
        chicken_rice_dim[23][14] = 16'b01101_010110_00111;
        chicken_rice_dim[23][15] = 16'b01101_010110_00111;
        chicken_rice_dim[23][16] = 16'b01000_010001_00100;
        chicken_rice_dim[23][17] = 16'b01001_010010_00101;
        chicken_rice_dim[23][18] = 16'b01001_010010_00101;
        chicken_rice_dim[23][19] = 16'b01000_010001_00100;
        chicken_rice_dim[23][20] = 16'b00111_001111_00100;
        chicken_rice_dim[23][21] = 16'b01010_010011_00101;
        chicken_rice_dim[23][22] = 16'b01000_010001_00100;
        chicken_rice_dim[23][23] = 16'b01010_010011_00101;
        chicken_rice_dim[23][24] = 16'b00110_001110_00011;
        chicken_rice_dim[23][25] = 16'b00110_001101_00010;
        chicken_rice_dim[23][26] = 16'b01011_011011_01111;
        chicken_rice_dim[23][27] = 16'b01011_011011_01111;
        chicken_rice_dim[23][28] = 16'b01011_011011_01111;
        chicken_rice_dim[23][29] = 16'b01011_011011_01111;
        chicken_rice_dim[23][30] = 16'b01011_011011_01111;
        chicken_rice_dim[23][31] = 16'b01011_011011_01111;
        chicken_rice_dim[24][0] = 16'b01011_011011_01111;
        chicken_rice_dim[24][1] = 16'b01011_011011_01111;
        chicken_rice_dim[24][2] = 16'b01011_011011_01111;
        chicken_rice_dim[24][3] = 16'b01011_011011_01111;
        chicken_rice_dim[24][4] = 16'b01011_011011_01111;
        chicken_rice_dim[24][5] = 16'b01011_011011_01111;
        chicken_rice_dim[24][6] = 16'b01011_011011_01111;
        chicken_rice_dim[24][7] = 16'b01011_011011_01111;
        chicken_rice_dim[24][8] = 16'b01011_011011_01111;
        chicken_rice_dim[24][9] = 16'b01011_011011_01111;
        chicken_rice_dim[24][10] = 16'b01101_010111_00111;
        chicken_rice_dim[24][11] = 16'b01110_011000_01000;
        chicken_rice_dim[24][12] = 16'b01110_011000_01000;
        chicken_rice_dim[24][13] = 16'b01101_011000_01000;
        chicken_rice_dim[24][14] = 16'b01101_010111_00111;
        chicken_rice_dim[24][15] = 16'b01101_010111_00111;
        chicken_rice_dim[24][16] = 16'b01101_010110_00111;
        chicken_rice_dim[24][17] = 16'b00111_001110_00011;
        chicken_rice_dim[24][18] = 16'b01000_010000_00100;
        chicken_rice_dim[24][19] = 16'b01000_010000_00100;
        chicken_rice_dim[24][20] = 16'b01001_010010_00101;
        chicken_rice_dim[24][21] = 16'b01000_010001_00100;
        chicken_rice_dim[24][22] = 16'b01000_010000_00100;
        chicken_rice_dim[24][23] = 16'b01001_010001_00100;
        chicken_rice_dim[24][24] = 16'b00110_001101_00011;
        chicken_rice_dim[24][25] = 16'b01011_011011_01111;
        chicken_rice_dim[24][26] = 16'b01011_011011_01111;
        chicken_rice_dim[24][27] = 16'b01011_011011_01111;
        chicken_rice_dim[24][28] = 16'b01011_011011_01111;
        chicken_rice_dim[24][29] = 16'b01011_011011_01111;
        chicken_rice_dim[24][30] = 16'b01011_011011_01111;
        chicken_rice_dim[24][31] = 16'b01011_011011_01111;
        chicken_rice_dim[25][0] = 16'b01011_011011_01111;
        chicken_rice_dim[25][1] = 16'b01011_011011_01111;
        chicken_rice_dim[25][2] = 16'b01011_011011_01111;
        chicken_rice_dim[25][3] = 16'b01011_011011_01111;
        chicken_rice_dim[25][4] = 16'b01011_011011_01111;
        chicken_rice_dim[25][5] = 16'b01011_011011_01111;
        chicken_rice_dim[25][6] = 16'b01011_011011_01111;
        chicken_rice_dim[25][7] = 16'b01011_011011_01111;
        chicken_rice_dim[25][8] = 16'b01011_011011_01111;
        chicken_rice_dim[25][9] = 16'b01011_011011_01111;
        chicken_rice_dim[25][10] = 16'b01011_011011_01111;
        chicken_rice_dim[25][11] = 16'b01011_011011_01111;
        chicken_rice_dim[25][12] = 16'b01011_011011_01111;
        chicken_rice_dim[25][13] = 16'b01011_011011_01111;
        chicken_rice_dim[25][14] = 16'b01011_011011_01111;
        chicken_rice_dim[25][15] = 16'b01011_011011_01111;
        chicken_rice_dim[25][16] = 16'b01011_011011_01111;
        chicken_rice_dim[25][17] = 16'b01011_011011_01111;
        chicken_rice_dim[25][18] = 16'b00110_001100_00010;
        chicken_rice_dim[25][19] = 16'b01000_010000_00011;
        chicken_rice_dim[25][20] = 16'b01001_010010_00100;
        chicken_rice_dim[25][21] = 16'b01010_010100_00110;
        chicken_rice_dim[25][22] = 16'b00110_001101_00010;
        chicken_rice_dim[25][23] = 16'b00111_001111_00011;
        chicken_rice_dim[25][24] = 16'b01011_011011_01111;
        chicken_rice_dim[25][25] = 16'b01011_011011_01111;
        chicken_rice_dim[25][26] = 16'b01011_011011_01111;
        chicken_rice_dim[25][27] = 16'b01011_011011_01111;
        chicken_rice_dim[25][28] = 16'b01011_011011_01111;
        chicken_rice_dim[25][29] = 16'b01011_011011_01111;
        chicken_rice_dim[25][30] = 16'b01011_011011_01111;
        chicken_rice_dim[25][31] = 16'b01011_011011_01111;
        chicken_rice_dim[26][0] = 16'b01011_011011_01111;
        chicken_rice_dim[26][1] = 16'b01011_011011_01111;
        chicken_rice_dim[26][2] = 16'b01011_011011_01111;
        chicken_rice_dim[26][3] = 16'b01011_011011_01111;
        chicken_rice_dim[26][4] = 16'b01011_011011_01111;
        chicken_rice_dim[26][5] = 16'b01011_011011_01111;
        chicken_rice_dim[26][6] = 16'b01011_011011_01111;
        chicken_rice_dim[26][7] = 16'b01011_011011_01111;
        chicken_rice_dim[26][8] = 16'b01011_011011_01111;
        chicken_rice_dim[26][9] = 16'b01011_011011_01111;
        chicken_rice_dim[26][10] = 16'b01011_011011_01111;
        chicken_rice_dim[26][11] = 16'b01011_011011_01111;
        chicken_rice_dim[26][12] = 16'b01011_011011_01111;
        chicken_rice_dim[26][13] = 16'b01011_011011_01111;
        chicken_rice_dim[26][14] = 16'b01011_011011_01111;
        chicken_rice_dim[26][15] = 16'b01011_011011_01111;
        chicken_rice_dim[26][16] = 16'b01011_011011_01111;
        chicken_rice_dim[26][17] = 16'b01011_011011_01111;
        chicken_rice_dim[26][18] = 16'b01011_011011_01111;
        chicken_rice_dim[26][19] = 16'b00110_001100_00010;
        chicken_rice_dim[26][20] = 16'b00110_001101_00010;
        chicken_rice_dim[26][21] = 16'b00110_001101_00011;
        chicken_rice_dim[26][22] = 16'b00101_001011_00010;
        chicken_rice_dim[26][23] = 16'b01011_011011_01111;
        chicken_rice_dim[26][24] = 16'b01011_011011_01111;
        chicken_rice_dim[26][25] = 16'b01011_011011_01111;
        chicken_rice_dim[26][26] = 16'b01011_011011_01111;
        chicken_rice_dim[26][27] = 16'b01011_011011_01111;
        chicken_rice_dim[26][28] = 16'b01011_011011_01111;
        chicken_rice_dim[26][29] = 16'b01011_011011_01111;
        chicken_rice_dim[26][30] = 16'b01011_011011_01111;
        chicken_rice_dim[26][31] = 16'b01011_011011_01111;
        chicken_rice_dim[27][0] = 16'b01011_011011_01111;
        chicken_rice_dim[27][1] = 16'b01011_011011_01111;
        chicken_rice_dim[27][2] = 16'b01011_011011_01111;
        chicken_rice_dim[27][3] = 16'b01011_011011_01111;
        chicken_rice_dim[27][4] = 16'b01011_011011_01111;
        chicken_rice_dim[27][5] = 16'b01011_011011_01111;
        chicken_rice_dim[27][6] = 16'b01011_011011_01111;
        chicken_rice_dim[27][7] = 16'b01011_011011_01111;
        chicken_rice_dim[27][8] = 16'b01011_011011_01111;
        chicken_rice_dim[27][9] = 16'b01011_011011_01111;
        chicken_rice_dim[27][10] = 16'b01011_011011_01111;
        chicken_rice_dim[27][11] = 16'b01011_011011_01111;
        chicken_rice_dim[27][12] = 16'b01011_011011_01111;
        chicken_rice_dim[27][13] = 16'b01011_011011_01111;
        chicken_rice_dim[27][14] = 16'b01011_011011_01111;
        chicken_rice_dim[27][15] = 16'b01011_011011_01111;
        chicken_rice_dim[27][16] = 16'b01011_011011_01111;
        chicken_rice_dim[27][17] = 16'b01011_011011_01111;
        chicken_rice_dim[27][18] = 16'b01011_011011_01111;
        chicken_rice_dim[27][19] = 16'b01011_011011_01111;
        chicken_rice_dim[27][20] = 16'b01011_011011_01111;
        chicken_rice_dim[27][21] = 16'b01011_011011_01111;
        chicken_rice_dim[27][22] = 16'b01011_011011_01111;
        chicken_rice_dim[27][23] = 16'b01011_011011_01111;
        chicken_rice_dim[27][24] = 16'b01011_011011_01111;
        chicken_rice_dim[27][25] = 16'b01011_011011_01111;
        chicken_rice_dim[27][26] = 16'b01011_011011_01111;
        chicken_rice_dim[27][27] = 16'b01011_011011_01111;
        chicken_rice_dim[27][28] = 16'b01011_011011_01111;
        chicken_rice_dim[27][29] = 16'b01011_011011_01111;
        chicken_rice_dim[27][30] = 16'b01011_011011_01111;
        chicken_rice_dim[27][31] = 16'b01011_011011_01111;
        chicken_rice_dim[28][0] = 16'b01011_011011_01111;
        chicken_rice_dim[28][1] = 16'b01011_011011_01111;
        chicken_rice_dim[28][2] = 16'b01011_011011_01111;
        chicken_rice_dim[28][3] = 16'b01011_011011_01111;
        chicken_rice_dim[28][4] = 16'b01011_011011_01111;
        chicken_rice_dim[28][5] = 16'b01011_011011_01111;
        chicken_rice_dim[28][6] = 16'b01011_011011_01111;
        chicken_rice_dim[28][7] = 16'b01011_011011_01111;
        chicken_rice_dim[28][8] = 16'b01011_011011_01111;
        chicken_rice_dim[28][9] = 16'b01011_011011_01111;
        chicken_rice_dim[28][10] = 16'b01011_011011_01111;
        chicken_rice_dim[28][11] = 16'b01011_011011_01111;
        chicken_rice_dim[28][12] = 16'b01011_011011_01111;
        chicken_rice_dim[28][13] = 16'b01011_011011_01111;
        chicken_rice_dim[28][14] = 16'b01011_011011_01111;
        chicken_rice_dim[28][15] = 16'b01011_011011_01111;
        chicken_rice_dim[28][16] = 16'b01011_011011_01111;
        chicken_rice_dim[28][17] = 16'b01011_011011_01111;
        chicken_rice_dim[28][18] = 16'b01011_011011_01111;
        chicken_rice_dim[28][19] = 16'b01011_011011_01111;
        chicken_rice_dim[28][20] = 16'b01011_011011_01111;
        chicken_rice_dim[28][21] = 16'b01011_011011_01111;
        chicken_rice_dim[28][22] = 16'b01011_011011_01111;
        chicken_rice_dim[28][23] = 16'b01011_011011_01111;
        chicken_rice_dim[28][24] = 16'b01011_011011_01111;
        chicken_rice_dim[28][25] = 16'b01011_011011_01111;
        chicken_rice_dim[28][26] = 16'b01011_011011_01111;
        chicken_rice_dim[28][27] = 16'b01011_011011_01111;
        chicken_rice_dim[28][28] = 16'b01011_011011_01111;
        chicken_rice_dim[28][29] = 16'b01011_011011_01111;
        chicken_rice_dim[28][30] = 16'b01011_011011_01111;
        chicken_rice_dim[28][31] = 16'b01011_011011_01111;
        chicken_rice_dim[29][0] = 16'b01011_011011_01111;
        chicken_rice_dim[29][1] = 16'b01011_011011_01111;
        chicken_rice_dim[29][2] = 16'b01011_011011_01111;
        chicken_rice_dim[29][3] = 16'b01011_011011_01111;
        chicken_rice_dim[29][4] = 16'b01011_011011_01111;
        chicken_rice_dim[29][5] = 16'b01011_011011_01111;
        chicken_rice_dim[29][6] = 16'b01011_011011_01111;
        chicken_rice_dim[29][7] = 16'b01011_011011_01111;
        chicken_rice_dim[29][8] = 16'b01011_011011_01111;
        chicken_rice_dim[29][9] = 16'b01011_011011_01111;
        chicken_rice_dim[29][10] = 16'b01011_011011_01111;
        chicken_rice_dim[29][11] = 16'b01011_011011_01111;
        chicken_rice_dim[29][12] = 16'b01011_011011_01111;
        chicken_rice_dim[29][13] = 16'b01011_011011_01111;
        chicken_rice_dim[29][14] = 16'b01011_011011_01111;
        chicken_rice_dim[29][15] = 16'b01011_011011_01111;
        chicken_rice_dim[29][16] = 16'b01011_011011_01111;
        chicken_rice_dim[29][17] = 16'b01011_011011_01111;
        chicken_rice_dim[29][18] = 16'b01011_011011_01111;
        chicken_rice_dim[29][19] = 16'b01011_011011_01111;
        chicken_rice_dim[29][20] = 16'b01011_011011_01111;
        chicken_rice_dim[29][21] = 16'b01011_011011_01111;
        chicken_rice_dim[29][22] = 16'b01011_011011_01111;
        chicken_rice_dim[29][23] = 16'b01011_011011_01111;
        chicken_rice_dim[29][24] = 16'b01011_011011_01111;
        chicken_rice_dim[29][25] = 16'b01011_011011_01111;
        chicken_rice_dim[29][26] = 16'b01011_011011_01111;
        chicken_rice_dim[29][27] = 16'b01011_011011_01111;
        chicken_rice_dim[29][28] = 16'b01011_011011_01111;
        chicken_rice_dim[29][29] = 16'b01011_011011_01111;
        chicken_rice_dim[29][30] = 16'b01011_011011_01111;
        chicken_rice_dim[29][31] = 16'b01011_011011_01111;
        chicken_rice_dim[30][0] = 16'b01011_011011_01111;
        chicken_rice_dim[30][1] = 16'b01011_011011_01111;
        chicken_rice_dim[30][2] = 16'b01011_011011_01111;
        chicken_rice_dim[30][3] = 16'b01011_011011_01111;
        chicken_rice_dim[30][4] = 16'b01011_011011_01111;
        chicken_rice_dim[30][5] = 16'b01011_011011_01111;
        chicken_rice_dim[30][6] = 16'b01011_011011_01111;
        chicken_rice_dim[30][7] = 16'b01011_011011_01111;
        chicken_rice_dim[30][8] = 16'b01011_011011_01111;
        chicken_rice_dim[30][9] = 16'b01011_011011_01111;
        chicken_rice_dim[30][10] = 16'b01011_011011_01111;
        chicken_rice_dim[30][11] = 16'b01011_011011_01111;
        chicken_rice_dim[30][12] = 16'b01011_011011_01111;
        chicken_rice_dim[30][13] = 16'b01011_011011_01111;
        chicken_rice_dim[30][14] = 16'b01011_011011_01111;
        chicken_rice_dim[30][15] = 16'b01011_011011_01111;
        chicken_rice_dim[30][16] = 16'b01011_011011_01111;
        chicken_rice_dim[30][17] = 16'b01011_011011_01111;
        chicken_rice_dim[30][18] = 16'b01011_011011_01111;
        chicken_rice_dim[30][19] = 16'b01011_011011_01111;
        chicken_rice_dim[30][20] = 16'b01011_011011_01111;
        chicken_rice_dim[30][21] = 16'b01011_011011_01111;
        chicken_rice_dim[30][22] = 16'b01011_011011_01111;
        chicken_rice_dim[30][23] = 16'b01011_011011_01111;
        chicken_rice_dim[30][24] = 16'b01011_011011_01111;
        chicken_rice_dim[30][25] = 16'b01011_011011_01111;
        chicken_rice_dim[30][26] = 16'b01011_011011_01111;
        chicken_rice_dim[30][27] = 16'b01011_011011_01111;
        chicken_rice_dim[30][28] = 16'b01011_011011_01111;
        chicken_rice_dim[30][29] = 16'b01011_011011_01111;
        chicken_rice_dim[30][30] = 16'b01011_011011_01111;
        chicken_rice_dim[30][31] = 16'b01011_011011_01111;
        chicken_rice_dim[31][0] = 16'b01011_011011_01111;
        chicken_rice_dim[31][1] = 16'b01011_011011_01111;
        chicken_rice_dim[31][2] = 16'b01011_011011_01111;
        chicken_rice_dim[31][3] = 16'b01011_011011_01111;
        chicken_rice_dim[31][4] = 16'b01011_011011_01111;
        chicken_rice_dim[31][5] = 16'b01011_011011_01111;
        chicken_rice_dim[31][6] = 16'b01011_011011_01111;
        chicken_rice_dim[31][7] = 16'b01011_011011_01111;
        chicken_rice_dim[31][8] = 16'b01011_011011_01111;
        chicken_rice_dim[31][9] = 16'b01011_011011_01111;
        chicken_rice_dim[31][10] = 16'b01011_011011_01111;
        chicken_rice_dim[31][11] = 16'b01011_011011_01111;
        chicken_rice_dim[31][12] = 16'b01011_011011_01111;
        chicken_rice_dim[31][13] = 16'b01011_011011_01111;
        chicken_rice_dim[31][14] = 16'b01011_011011_01111;
        chicken_rice_dim[31][15] = 16'b01011_011011_01111;
        chicken_rice_dim[31][16] = 16'b01011_011011_01111;
        chicken_rice_dim[31][17] = 16'b01011_011011_01111;
        chicken_rice_dim[31][18] = 16'b01011_011011_01111;
        chicken_rice_dim[31][19] = 16'b01011_011011_01111;
        chicken_rice_dim[31][20] = 16'b01011_011011_01111;
        chicken_rice_dim[31][21] = 16'b01011_011011_01111;
        chicken_rice_dim[31][22] = 16'b01011_011011_01111;
        chicken_rice_dim[31][23] = 16'b01011_011011_01111;
        chicken_rice_dim[31][24] = 16'b01011_011011_01111;
        chicken_rice_dim[31][25] = 16'b01011_011011_01111;
        chicken_rice_dim[31][26] = 16'b01011_011011_01111;
        chicken_rice_dim[31][27] = 16'b01011_011011_01111;
        chicken_rice_dim[31][28] = 16'b01011_011011_01111;
        chicken_rice_dim[31][29] = 16'b01011_011011_01111;
        chicken_rice_dim[31][30] = 16'b01011_011011_01111;
        chicken_rice_dim[31][31] = 16'b01011_011011_01111;
        
        
                
        onion_soup_dim[0][0] = 16'b01111_010101_01010;
        onion_soup_dim[0][1] = 16'b01111_010101_01010;
        onion_soup_dim[0][2] = 16'b01111_010101_01010;
        onion_soup_dim[0][3] = 16'b01111_010101_01010;
        onion_soup_dim[0][4] = 16'b01111_010101_01010;
        onion_soup_dim[0][5] = 16'b01111_010101_01010;
        onion_soup_dim[0][6] = 16'b01111_010101_01010;
        onion_soup_dim[0][7] = 16'b01111_010101_01010;
        onion_soup_dim[0][8] = 16'b01111_010101_01010;
        onion_soup_dim[0][9] = 16'b01111_010101_01010;
        onion_soup_dim[0][10] = 16'b01111_010101_01010;
        onion_soup_dim[0][11] = 16'b01111_010101_01010;
        onion_soup_dim[0][12] = 16'b01111_010101_01010;
        onion_soup_dim[0][13] = 16'b01111_010101_01010;
        onion_soup_dim[0][14] = 16'b01111_010101_01010;
        onion_soup_dim[0][15] = 16'b01111_010101_01010;
        onion_soup_dim[0][16] = 16'b01111_010101_01010;
        onion_soup_dim[0][17] = 16'b01111_010101_01010;
        onion_soup_dim[0][18] = 16'b01111_010101_01010;
        onion_soup_dim[0][19] = 16'b01111_010101_01010;
        onion_soup_dim[0][20] = 16'b01111_010101_01010;
        onion_soup_dim[0][21] = 16'b01111_010101_01010;
        onion_soup_dim[0][22] = 16'b01111_010101_01010;
        onion_soup_dim[0][23] = 16'b01111_010101_01010;
        onion_soup_dim[0][24] = 16'b01111_010101_01010;
        onion_soup_dim[0][25] = 16'b01111_010101_01010;
        onion_soup_dim[0][26] = 16'b01111_010101_01010;
        onion_soup_dim[0][27] = 16'b01111_010101_01010;
        onion_soup_dim[0][28] = 16'b01111_010101_01010;
        onion_soup_dim[0][29] = 16'b01111_010101_01010;
        onion_soup_dim[0][30] = 16'b01111_010101_01010;
        onion_soup_dim[0][31] = 16'b01111_010101_01010;
        onion_soup_dim[1][0] = 16'b01111_010101_01010;
        onion_soup_dim[1][1] = 16'b01111_010101_01010;
        onion_soup_dim[1][2] = 16'b01111_010101_01010;
        onion_soup_dim[1][3] = 16'b01111_010101_01010;
        onion_soup_dim[1][4] = 16'b01111_010101_01010;
        onion_soup_dim[1][5] = 16'b01111_010101_01010;
        onion_soup_dim[1][6] = 16'b01111_010101_01010;
        onion_soup_dim[1][7] = 16'b01111_010101_01010;
        onion_soup_dim[1][8] = 16'b01111_010101_01010;
        onion_soup_dim[1][9] = 16'b01111_010101_01010;
        onion_soup_dim[1][10] = 16'b01111_010101_01010;
        onion_soup_dim[1][11] = 16'b01111_010101_01010;
        onion_soup_dim[1][12] = 16'b01111_010101_01010;
        onion_soup_dim[1][13] = 16'b01111_010101_01010;
        onion_soup_dim[1][14] = 16'b01111_010101_01010;
        onion_soup_dim[1][15] = 16'b01111_010101_01010;
        onion_soup_dim[1][16] = 16'b01111_010101_01010;
        onion_soup_dim[1][17] = 16'b01111_010101_01010;
        onion_soup_dim[1][18] = 16'b01111_010101_01010;
        onion_soup_dim[1][19] = 16'b01111_010101_01010;
        onion_soup_dim[1][20] = 16'b01111_010101_01010;
        onion_soup_dim[1][21] = 16'b01111_010101_01010;
        onion_soup_dim[1][22] = 16'b01111_010101_01010;
        onion_soup_dim[1][23] = 16'b01111_010101_01010;
        onion_soup_dim[1][24] = 16'b01111_010101_01010;
        onion_soup_dim[1][25] = 16'b01111_010101_01010;
        onion_soup_dim[1][26] = 16'b01111_010101_01010;
        onion_soup_dim[1][27] = 16'b01111_010101_01010;
        onion_soup_dim[1][28] = 16'b01111_010101_01010;
        onion_soup_dim[1][29] = 16'b01111_010101_01010;
        onion_soup_dim[1][30] = 16'b01111_010101_01010;
        onion_soup_dim[1][31] = 16'b01111_010101_01010;
        onion_soup_dim[2][0] = 16'b01111_010101_01010;
        onion_soup_dim[2][1] = 16'b01111_010101_01010;
        onion_soup_dim[2][2] = 16'b01111_010101_01010;
        onion_soup_dim[2][3] = 16'b01111_010101_01010;
        onion_soup_dim[2][4] = 16'b01111_010101_01010;
        onion_soup_dim[2][5] = 16'b01111_010101_01010;
        onion_soup_dim[2][6] = 16'b01111_010101_01010;
        onion_soup_dim[2][7] = 16'b01111_010101_01010;
        onion_soup_dim[2][8] = 16'b01111_010101_01010;
        onion_soup_dim[2][9] = 16'b01111_010101_01010;
        onion_soup_dim[2][10] = 16'b01111_010101_01010;
        onion_soup_dim[2][11] = 16'b01111_010101_01010;
        onion_soup_dim[2][12] = 16'b01111_010101_01010;
        onion_soup_dim[2][13] = 16'b01111_010101_01010;
        onion_soup_dim[2][14] = 16'b01111_010101_01010;
        onion_soup_dim[2][15] = 16'b01111_010101_01010;
        onion_soup_dim[2][16] = 16'b01111_010101_01010;
        onion_soup_dim[2][17] = 16'b01111_010101_01010;
        onion_soup_dim[2][18] = 16'b01111_010101_01010;
        onion_soup_dim[2][19] = 16'b01111_010101_01010;
        onion_soup_dim[2][20] = 16'b01111_010101_01010;
        onion_soup_dim[2][21] = 16'b01111_010101_01010;
        onion_soup_dim[2][22] = 16'b01111_010101_01010;
        onion_soup_dim[2][23] = 16'b01111_010101_01010;
        onion_soup_dim[2][24] = 16'b01111_010101_01010;
        onion_soup_dim[2][25] = 16'b01111_010101_01010;
        onion_soup_dim[2][26] = 16'b01111_010101_01010;
        onion_soup_dim[2][27] = 16'b01111_010101_01010;
        onion_soup_dim[2][28] = 16'b01111_010101_01010;
        onion_soup_dim[2][29] = 16'b01111_010101_01010;
        onion_soup_dim[2][30] = 16'b01111_010101_01010;
        onion_soup_dim[2][31] = 16'b01111_010101_01010;
        onion_soup_dim[3][0] = 16'b01111_010101_01010;
        onion_soup_dim[3][1] = 16'b01111_010101_01010;
        onion_soup_dim[3][2] = 16'b01111_010101_01010;
        onion_soup_dim[3][3] = 16'b01111_010101_01010;
        onion_soup_dim[3][4] = 16'b01111_010101_01010;
        onion_soup_dim[3][5] = 16'b01111_010101_01010;
        onion_soup_dim[3][6] = 16'b01111_010101_01010;
        onion_soup_dim[3][7] = 16'b01111_010101_01010;
        onion_soup_dim[3][8] = 16'b01111_010101_01010;
        onion_soup_dim[3][9] = 16'b01111_010101_01010;
        onion_soup_dim[3][10] = 16'b01111_010101_01010;
        onion_soup_dim[3][11] = 16'b01111_010101_01010;
        onion_soup_dim[3][12] = 16'b01111_010101_01010;
        onion_soup_dim[3][13] = 16'b01111_010101_01010;
        onion_soup_dim[3][14] = 16'b01111_010101_01010;
        onion_soup_dim[3][15] = 16'b01111_010101_01010;
        onion_soup_dim[3][16] = 16'b01111_010101_01010;
        onion_soup_dim[3][17] = 16'b01111_010101_01010;
        onion_soup_dim[3][18] = 16'b01111_010101_01010;
        onion_soup_dim[3][19] = 16'b01111_010101_01010;
        onion_soup_dim[3][20] = 16'b01111_010101_01010;
        onion_soup_dim[3][21] = 16'b01111_010101_01010;
        onion_soup_dim[3][22] = 16'b01111_010101_01010;
        onion_soup_dim[3][23] = 16'b01111_010101_01010;
        onion_soup_dim[3][24] = 16'b01111_010101_01010;
        onion_soup_dim[3][25] = 16'b01111_010101_01010;
        onion_soup_dim[3][26] = 16'b01111_010101_01010;
        onion_soup_dim[3][27] = 16'b01111_010101_01010;
        onion_soup_dim[3][28] = 16'b01111_010101_01010;
        onion_soup_dim[3][29] = 16'b01111_010101_01010;
        onion_soup_dim[3][30] = 16'b01111_010101_01010;
        onion_soup_dim[3][31] = 16'b01111_010101_01010;
        onion_soup_dim[4][0] = 16'b01111_010101_01010;
        onion_soup_dim[4][1] = 16'b01111_010101_01010;
        onion_soup_dim[4][2] = 16'b01111_010101_01010;
        onion_soup_dim[4][3] = 16'b01111_010101_01010;
        onion_soup_dim[4][4] = 16'b01111_010101_01010;
        onion_soup_dim[4][5] = 16'b01111_010101_01010;
        onion_soup_dim[4][6] = 16'b01111_010101_01010;
        onion_soup_dim[4][7] = 16'b01111_010101_01010;
        onion_soup_dim[4][8] = 16'b01111_010101_01010;
        onion_soup_dim[4][9] = 16'b01111_010101_01010;
        onion_soup_dim[4][10] = 16'b01111_010101_01010;
        onion_soup_dim[4][11] = 16'b01111_010101_01010;
        onion_soup_dim[4][12] = 16'b01111_010101_01010;
        onion_soup_dim[4][13] = 16'b01111_010101_01010;
        onion_soup_dim[4][14] = 16'b01111_010101_01010;
        onion_soup_dim[4][15] = 16'b01111_010101_01010;
        onion_soup_dim[4][16] = 16'b01111_010101_01010;
        onion_soup_dim[4][17] = 16'b01111_010101_01010;
        onion_soup_dim[4][18] = 16'b01111_010101_01010;
        onion_soup_dim[4][19] = 16'b01111_010101_01010;
        onion_soup_dim[4][20] = 16'b01111_010101_01010;
        onion_soup_dim[4][21] = 16'b01111_010101_01010;
        onion_soup_dim[4][22] = 16'b01111_010101_01010;
        onion_soup_dim[4][23] = 16'b01111_010101_01010;
        onion_soup_dim[4][24] = 16'b01111_010101_01010;
        onion_soup_dim[4][25] = 16'b01111_010101_01010;
        onion_soup_dim[4][26] = 16'b01111_010101_01010;
        onion_soup_dim[4][27] = 16'b01111_010101_01010;
        onion_soup_dim[4][28] = 16'b01111_010101_01010;
        onion_soup_dim[4][29] = 16'b01111_010101_01010;
        onion_soup_dim[4][30] = 16'b01111_010101_01010;
        onion_soup_dim[4][31] = 16'b01111_010101_01010;
        onion_soup_dim[5][0] = 16'b01111_010101_01010;
        onion_soup_dim[5][1] = 16'b01111_010101_01010;
        onion_soup_dim[5][2] = 16'b01111_010101_01010;
        onion_soup_dim[5][3] = 16'b01111_010101_01010;
        onion_soup_dim[5][4] = 16'b01111_010101_01010;
        onion_soup_dim[5][5] = 16'b01111_010101_01010;
        onion_soup_dim[5][6] = 16'b01111_010101_01010;
        onion_soup_dim[5][7] = 16'b01111_010101_01010;
        onion_soup_dim[5][8] = 16'b01111_010101_01010;
        onion_soup_dim[5][9] = 16'b01111_010101_01010;
        onion_soup_dim[5][10] = 16'b01111_010101_01010;
        onion_soup_dim[5][11] = 16'b01111_010101_01010;
        onion_soup_dim[5][12] = 16'b01111_010101_01010;
        onion_soup_dim[5][13] = 16'b01111_010101_01010;
        onion_soup_dim[5][14] = 16'b01111_010101_01010;
        onion_soup_dim[5][15] = 16'b01111_010101_01010;
        onion_soup_dim[5][16] = 16'b01111_010101_01010;
        onion_soup_dim[5][17] = 16'b01111_010101_01010;
        onion_soup_dim[5][18] = 16'b01111_010101_01010;
        onion_soup_dim[5][19] = 16'b01111_010101_01010;
        onion_soup_dim[5][20] = 16'b01111_010101_01010;
        onion_soup_dim[5][21] = 16'b01111_010101_01010;
        onion_soup_dim[5][22] = 16'b01111_010101_01010;
        onion_soup_dim[5][23] = 16'b01111_010101_01010;
        onion_soup_dim[5][24] = 16'b01111_010101_01010;
        onion_soup_dim[5][25] = 16'b01111_010101_01010;
        onion_soup_dim[5][26] = 16'b01111_010101_01010;
        onion_soup_dim[5][27] = 16'b01111_010101_01010;
        onion_soup_dim[5][28] = 16'b01111_010101_01010;
        onion_soup_dim[5][29] = 16'b01111_010101_01010;
        onion_soup_dim[5][30] = 16'b01111_010101_01010;
        onion_soup_dim[5][31] = 16'b01111_010101_01010;
        onion_soup_dim[6][0] = 16'b01111_010101_01010;
        onion_soup_dim[6][1] = 16'b01111_010101_01010;
        onion_soup_dim[6][2] = 16'b01111_010101_01010;
        onion_soup_dim[6][3] = 16'b01111_010101_01010;
        onion_soup_dim[6][4] = 16'b01111_010101_01010;
        onion_soup_dim[6][5] = 16'b01111_010101_01010;
        onion_soup_dim[6][6] = 16'b01111_010101_01010;
        onion_soup_dim[6][7] = 16'b01111_010101_01010;
        onion_soup_dim[6][8] = 16'b01111_010101_01010;
        onion_soup_dim[6][9] = 16'b01111_010101_01010;
        onion_soup_dim[6][10] = 16'b01111_010101_01010;
        onion_soup_dim[6][11] = 16'b01111_010101_01010;
        onion_soup_dim[6][12] = 16'b01000_001010_00001;
        onion_soup_dim[6][13] = 16'b01000_001010_00001;
        onion_soup_dim[6][14] = 16'b01010_001101_00010;
        onion_soup_dim[6][15] = 16'b01001_001011_00001;
        onion_soup_dim[6][16] = 16'b01001_001010_00001;
        onion_soup_dim[6][17] = 16'b01000_001010_00001;
        onion_soup_dim[6][18] = 16'b01001_001011_00001;
        onion_soup_dim[6][19] = 16'b01001_001100_00010;
        onion_soup_dim[6][20] = 16'b01000_001010_00001;
        onion_soup_dim[6][21] = 16'b01111_010101_01010;
        onion_soup_dim[6][22] = 16'b01111_010101_01010;
        onion_soup_dim[6][23] = 16'b01111_010101_01010;
        onion_soup_dim[6][24] = 16'b01111_010101_01010;
        onion_soup_dim[6][25] = 16'b01111_010101_01010;
        onion_soup_dim[6][26] = 16'b01111_010101_01010;
        onion_soup_dim[6][27] = 16'b01111_010101_01010;
        onion_soup_dim[6][28] = 16'b01111_010101_01010;
        onion_soup_dim[6][29] = 16'b01111_010101_01010;
        onion_soup_dim[6][30] = 16'b01111_010101_01010;
        onion_soup_dim[6][31] = 16'b01111_010101_01010;
        onion_soup_dim[7][0] = 16'b01111_010101_01010;
        onion_soup_dim[7][1] = 16'b01111_010101_01010;
        onion_soup_dim[7][2] = 16'b01111_010101_01010;
        onion_soup_dim[7][3] = 16'b01111_010101_01010;
        onion_soup_dim[7][4] = 16'b01111_010101_01010;
        onion_soup_dim[7][5] = 16'b01111_010101_01010;
        onion_soup_dim[7][6] = 16'b01111_010101_01010;
        onion_soup_dim[7][7] = 16'b01111_010101_01010;
        onion_soup_dim[7][8] = 16'b01111_010101_01010;
        onion_soup_dim[7][9] = 16'b01111_010101_01010;
        onion_soup_dim[7][10] = 16'b01000_001001_00001;
        onion_soup_dim[7][11] = 16'b00111_001001_00001;
        onion_soup_dim[7][12] = 16'b01001_001101_00010;
        onion_soup_dim[7][13] = 16'b01000_001011_00001;
        onion_soup_dim[7][14] = 16'b01011_001111_00011;
        onion_soup_dim[7][15] = 16'b01001_001011_00001;
        onion_soup_dim[7][16] = 16'b01011_001110_00011;
        onion_soup_dim[7][17] = 16'b01100_010001_00100;
        onion_soup_dim[7][18] = 16'b00111_001001_00001;
        onion_soup_dim[7][19] = 16'b01001_001100_00010;
        onion_soup_dim[7][20] = 16'b00111_001001_00001;
        onion_soup_dim[7][21] = 16'b01000_001001_00001;
        onion_soup_dim[7][22] = 16'b01000_001001_00001;
        onion_soup_dim[7][23] = 16'b01111_010101_01010;
        onion_soup_dim[7][24] = 16'b01111_010101_01010;
        onion_soup_dim[7][25] = 16'b01111_010101_01010;
        onion_soup_dim[7][26] = 16'b01111_010101_01010;
        onion_soup_dim[7][27] = 16'b01111_010101_01010;
        onion_soup_dim[7][28] = 16'b01111_010101_01010;
        onion_soup_dim[7][29] = 16'b01111_010101_01010;
        onion_soup_dim[7][30] = 16'b01111_010101_01010;
        onion_soup_dim[7][31] = 16'b01111_010101_01010;
        onion_soup_dim[8][0] = 16'b01111_010101_01010;
        onion_soup_dim[8][1] = 16'b01111_010101_01010;
        onion_soup_dim[8][2] = 16'b01111_010101_01010;
        onion_soup_dim[8][3] = 16'b01111_010101_01010;
        onion_soup_dim[8][4] = 16'b01111_010101_01010;
        onion_soup_dim[8][5] = 16'b01111_010101_01010;
        onion_soup_dim[8][6] = 16'b01111_010101_01010;
        onion_soup_dim[8][7] = 16'b01111_010101_01010;
        onion_soup_dim[8][8] = 16'b01010_001100_00010;
        onion_soup_dim[8][9] = 16'b01001_001100_00010;
        onion_soup_dim[8][10] = 16'b01011_010000_00011;
        onion_soup_dim[8][11] = 16'b01010_001101_00010;
        onion_soup_dim[8][12] = 16'b01010_001101_00010;
        onion_soup_dim[8][13] = 16'b01001_001100_00010;
        onion_soup_dim[8][14] = 16'b01001_001100_00010;
        onion_soup_dim[8][15] = 16'b01101_010011_00100;
        onion_soup_dim[8][16] = 16'b01010_001101_00010;
        onion_soup_dim[8][17] = 16'b01011_001110_00010;
        onion_soup_dim[8][18] = 16'b01001_001011_00010;
        onion_soup_dim[8][19] = 16'b01011_001111_00011;
        onion_soup_dim[8][20] = 16'b01000_001001_00001;
        onion_soup_dim[8][21] = 16'b01010_001101_00010;
        onion_soup_dim[8][22] = 16'b01010_001101_00010;
        onion_soup_dim[8][23] = 16'b01000_001001_00001;
        onion_soup_dim[8][24] = 16'b01111_010101_01010;
        onion_soup_dim[8][25] = 16'b01111_010101_01010;
        onion_soup_dim[8][26] = 16'b01111_010101_01010;
        onion_soup_dim[8][27] = 16'b01111_010101_01010;
        onion_soup_dim[8][28] = 16'b01111_010101_01010;
        onion_soup_dim[8][29] = 16'b01111_010101_01010;
        onion_soup_dim[8][30] = 16'b01111_010101_01010;
        onion_soup_dim[8][31] = 16'b01111_010101_01010;
        onion_soup_dim[9][0] = 16'b01111_010101_01010;
        onion_soup_dim[9][1] = 16'b01111_010101_01010;
        onion_soup_dim[9][2] = 16'b01111_010101_01010;
        onion_soup_dim[9][3] = 16'b01111_010101_01010;
        onion_soup_dim[9][4] = 16'b01111_010101_01010;
        onion_soup_dim[9][5] = 16'b01111_010101_01010;
        onion_soup_dim[9][6] = 16'b01111_010101_01010;
        onion_soup_dim[9][7] = 16'b01000_001010_00001;
        onion_soup_dim[9][8] = 16'b01010_001101_00010;
        onion_soup_dim[9][9] = 16'b01100_010010_00100;
        onion_soup_dim[9][10] = 16'b01100_010010_00100;
        onion_soup_dim[9][11] = 16'b01010_001110_00011;
        onion_soup_dim[9][12] = 16'b01011_001110_00011;
        onion_soup_dim[9][13] = 16'b01010_001101_00010;
        onion_soup_dim[9][14] = 16'b01101_010011_00100;
        onion_soup_dim[9][15] = 16'b01010_001101_00010;
        onion_soup_dim[9][16] = 16'b01001_001011_00001;
        onion_soup_dim[9][17] = 16'b01011_001111_00011;
        onion_soup_dim[9][18] = 16'b01011_001110_00010;
        onion_soup_dim[9][19] = 16'b01010_001110_00011;
        onion_soup_dim[9][20] = 16'b00111_000111_00001;
        onion_soup_dim[9][21] = 16'b01010_001101_00010;
        onion_soup_dim[9][22] = 16'b01011_001110_00011;
        onion_soup_dim[9][23] = 16'b01010_001100_00010;
        onion_soup_dim[9][24] = 16'b01001_001100_00010;
        onion_soup_dim[9][25] = 16'b01111_010101_01010;
        onion_soup_dim[9][26] = 16'b01111_010101_01010;
        onion_soup_dim[9][27] = 16'b01111_010101_01010;
        onion_soup_dim[9][28] = 16'b01111_010101_01010;
        onion_soup_dim[9][29] = 16'b01111_010101_01010;
        onion_soup_dim[9][30] = 16'b01111_010101_01010;
        onion_soup_dim[9][31] = 16'b01111_010101_01010;
        onion_soup_dim[10][0] = 16'b01111_010101_01010;
        onion_soup_dim[10][1] = 16'b01111_010101_01010;
        onion_soup_dim[10][2] = 16'b01111_010101_01010;
        onion_soup_dim[10][3] = 16'b01111_010101_01010;
        onion_soup_dim[10][4] = 16'b01111_010101_01010;
        onion_soup_dim[10][5] = 16'b01111_010101_01010;
        onion_soup_dim[10][6] = 16'b00110_000110_00000;
        onion_soup_dim[10][7] = 16'b01001_001011_00010;
        onion_soup_dim[10][8] = 16'b01010_001110_00010;
        onion_soup_dim[10][9] = 16'b01011_001110_00011;
        onion_soup_dim[10][10] = 16'b01101_010101_00101;
        onion_soup_dim[10][11] = 16'b01011_001111_00011;
        onion_soup_dim[10][12] = 16'b00110_000110_00000;
        onion_soup_dim[10][13] = 16'b01000_001001_00001;
        onion_soup_dim[10][14] = 16'b00101_000101_00000;
        onion_soup_dim[10][15] = 16'b00111_001000_00001;
        onion_soup_dim[10][16] = 16'b00110_000110_00000;
        onion_soup_dim[10][17] = 16'b01001_001011_00001;
        onion_soup_dim[10][18] = 16'b00111_001000_00000;
        onion_soup_dim[10][19] = 16'b01000_001001_00001;
        onion_soup_dim[10][20] = 16'b01000_001001_00001;
        onion_soup_dim[10][21] = 16'b00111_001001_00001;
        onion_soup_dim[10][22] = 16'b01010_001110_00010;
        onion_soup_dim[10][23] = 16'b01011_010000_00011;
        onion_soup_dim[10][24] = 16'b01000_001010_00001;
        onion_soup_dim[10][25] = 16'b01001_001011_00001;
        onion_soup_dim[10][26] = 16'b01000_001011_00001;
        onion_soup_dim[10][27] = 16'b01111_010101_01010;
        onion_soup_dim[10][28] = 16'b01111_010101_01010;
        onion_soup_dim[10][29] = 16'b01111_010101_01010;
        onion_soup_dim[10][30] = 16'b01111_010101_01010;
        onion_soup_dim[10][31] = 16'b01111_010101_01010;
        onion_soup_dim[11][0] = 16'b01111_010101_01010;
        onion_soup_dim[11][1] = 16'b01111_010101_01010;
        onion_soup_dim[11][2] = 16'b01111_010101_01010;
        onion_soup_dim[11][3] = 16'b01111_010101_01010;
        onion_soup_dim[11][4] = 16'b01111_010101_01010;
        onion_soup_dim[11][5] = 16'b01000_001010_00001;
        onion_soup_dim[11][6] = 16'b01010_001101_00010;
        onion_soup_dim[11][7] = 16'b01011_001110_00011;
        onion_soup_dim[11][8] = 16'b01010_001101_00010;
        onion_soup_dim[11][9] = 16'b00110_000111_00000;
        onion_soup_dim[11][10] = 16'b01001_001011_00001;
        onion_soup_dim[11][11] = 16'b01001_001011_00001;
        onion_soup_dim[11][12] = 16'b01000_001010_00001;
        onion_soup_dim[11][13] = 16'b01000_001001_00001;
        onion_soup_dim[11][14] = 16'b01001_001100_00001;
        onion_soup_dim[11][15] = 16'b01010_001100_00001;
        onion_soup_dim[11][16] = 16'b01001_001010_00001;
        onion_soup_dim[11][17] = 16'b01000_001010_00001;
        onion_soup_dim[11][18] = 16'b01000_001001_00001;
        onion_soup_dim[11][19] = 16'b01000_001001_00001;
        onion_soup_dim[11][20] = 16'b00111_001000_00001;
        onion_soup_dim[11][21] = 16'b00111_001000_00001;
        onion_soup_dim[11][22] = 16'b01000_001001_00001;
        onion_soup_dim[11][23] = 16'b00110_000111_00000;
        onion_soup_dim[11][24] = 16'b01010_001100_00010;
        onion_soup_dim[11][25] = 16'b01001_001100_00010;
        onion_soup_dim[11][26] = 16'b00111_001001_00001;
        onion_soup_dim[11][27] = 16'b01111_010101_01010;
        onion_soup_dim[11][28] = 16'b01111_010101_01010;
        onion_soup_dim[11][29] = 16'b01111_010101_01010;
        onion_soup_dim[11][30] = 16'b01111_010101_01010;
        onion_soup_dim[11][31] = 16'b01111_010101_01010;
        onion_soup_dim[12][0] = 16'b01111_010101_01010;
        onion_soup_dim[12][1] = 16'b01111_010101_01010;
        onion_soup_dim[12][2] = 16'b01111_010101_01010;
        onion_soup_dim[12][3] = 16'b01111_010101_01010;
        onion_soup_dim[12][4] = 16'b01111_010101_01010;
        onion_soup_dim[12][5] = 16'b01001_001101_00010;
        onion_soup_dim[12][6] = 16'b01010_001101_00010;
        onion_soup_dim[12][7] = 16'b00110_000111_00000;
        onion_soup_dim[12][8] = 16'b00111_001000_00001;
        onion_soup_dim[12][9] = 16'b00110_000110_00000;
        onion_soup_dim[12][10] = 16'b00110_000111_00000;
        onion_soup_dim[12][11] = 16'b00111_001000_00001;
        onion_soup_dim[12][12] = 16'b00101_000100_00000;
        onion_soup_dim[12][13] = 16'b00100_000100_00000;
        onion_soup_dim[12][14] = 16'b00110_000110_00000;
        onion_soup_dim[12][15] = 16'b00100_000011_00000;
        onion_soup_dim[12][16] = 16'b00111_001000_00000;
        onion_soup_dim[12][17] = 16'b00011_000011_00000;
        onion_soup_dim[12][18] = 16'b00101_000101_00000;
        onion_soup_dim[12][19] = 16'b00110_000110_00000;
        onion_soup_dim[12][20] = 16'b00110_000111_00000;
        onion_soup_dim[12][21] = 16'b01001_001010_00001;
        onion_soup_dim[12][22] = 16'b00111_001000_00001;
        onion_soup_dim[12][23] = 16'b01001_001011_00001;
        onion_soup_dim[12][24] = 16'b00101_000101_00000;
        onion_soup_dim[12][25] = 16'b01001_001100_00010;
        onion_soup_dim[12][26] = 16'b00100_000100_00000;
        onion_soup_dim[12][27] = 16'b01111_010101_01010;
        onion_soup_dim[12][28] = 16'b01111_010101_01010;
        onion_soup_dim[12][29] = 16'b01111_010101_01010;
        onion_soup_dim[12][30] = 16'b01111_010101_01010;
        onion_soup_dim[12][31] = 16'b01111_010101_01010;
        onion_soup_dim[13][0] = 16'b01111_010101_01010;
        onion_soup_dim[13][1] = 16'b01111_010101_01010;
        onion_soup_dim[13][2] = 16'b01111_010101_01010;
        onion_soup_dim[13][3] = 16'b01111_010101_01010;
        onion_soup_dim[13][4] = 16'b01100_010000_00011;
        onion_soup_dim[13][5] = 16'b00110_000111_00000;
        onion_soup_dim[13][6] = 16'b00111_001000_00001;
        onion_soup_dim[13][7] = 16'b01010_001101_00010;
        onion_soup_dim[13][8] = 16'b00110_000110_00000;
        onion_soup_dim[13][9] = 16'b00100_000100_00000;
        onion_soup_dim[13][10] = 16'b00101_000101_00000;
        onion_soup_dim[13][11] = 16'b00100_000100_00000;
        onion_soup_dim[13][12] = 16'b00101_000101_00000;
        onion_soup_dim[13][13] = 16'b01001_001011_00001;
        onion_soup_dim[13][14] = 16'b00100_000100_00000;
        onion_soup_dim[13][15] = 16'b00101_000101_00000;
        onion_soup_dim[13][16] = 16'b00111_001000_00001;
        onion_soup_dim[13][17] = 16'b00110_000111_00000;
        onion_soup_dim[13][18] = 16'b00110_000111_00000;
        onion_soup_dim[13][19] = 16'b00110_000111_00000;
        onion_soup_dim[13][20] = 16'b00101_000101_00000;
        onion_soup_dim[13][21] = 16'b00111_000111_00000;
        onion_soup_dim[13][22] = 16'b00110_000111_00000;
        onion_soup_dim[13][23] = 16'b00110_000110_00000;
        onion_soup_dim[13][24] = 16'b01000_001010_00001;
        onion_soup_dim[13][25] = 16'b01000_001001_00001;
        onion_soup_dim[13][26] = 16'b00111_001001_00001;
        onion_soup_dim[13][27] = 16'b01001_001011_00001;
        onion_soup_dim[13][28] = 16'b01111_010101_01010;
        onion_soup_dim[13][29] = 16'b01111_010101_01010;
        onion_soup_dim[13][30] = 16'b01111_010101_01010;
        onion_soup_dim[13][31] = 16'b01111_010101_01010;
        onion_soup_dim[14][0] = 16'b01111_010101_01010;
        onion_soup_dim[14][1] = 16'b01111_010101_01010;
        onion_soup_dim[14][2] = 16'b01111_010101_01010;
        onion_soup_dim[14][3] = 16'b01111_010101_01010;
        onion_soup_dim[14][4] = 16'b01001_001100_00010;
        onion_soup_dim[14][5] = 16'b00100_000100_00000;
        onion_soup_dim[14][6] = 16'b00111_001000_00000;
        onion_soup_dim[14][7] = 16'b00101_000110_00000;
        onion_soup_dim[14][8] = 16'b00101_000101_00000;
        onion_soup_dim[14][9] = 16'b00111_000111_00000;
        onion_soup_dim[14][10] = 16'b00110_000110_00000;
        onion_soup_dim[14][11] = 16'b00110_000110_00000;
        onion_soup_dim[14][12] = 16'b00101_000110_00000;
        onion_soup_dim[14][13] = 16'b00110_000110_00000;
        onion_soup_dim[14][14] = 16'b00100_000100_00000;
        onion_soup_dim[14][15] = 16'b00110_000110_00000;
        onion_soup_dim[14][16] = 16'b00100_000100_00000;
        onion_soup_dim[14][17] = 16'b01001_001101_00010;
        onion_soup_dim[14][18] = 16'b01011_001111_00011;
        onion_soup_dim[14][19] = 16'b00110_000111_00000;
        onion_soup_dim[14][20] = 16'b00110_000110_00000;
        onion_soup_dim[14][21] = 16'b00101_000110_00000;
        onion_soup_dim[14][22] = 16'b00110_000110_00000;
        onion_soup_dim[14][23] = 16'b00110_000110_00000;
        onion_soup_dim[14][24] = 16'b00101_000101_00000;
        onion_soup_dim[14][25] = 16'b00111_001000_00001;
        onion_soup_dim[14][26] = 16'b01000_001001_00001;
        onion_soup_dim[14][27] = 16'b01001_001100_00010;
        onion_soup_dim[14][28] = 16'b01111_010101_01010;
        onion_soup_dim[14][29] = 16'b01111_010101_01010;
        onion_soup_dim[14][30] = 16'b01111_010101_01010;
        onion_soup_dim[14][31] = 16'b01111_010101_01010;
        onion_soup_dim[15][0] = 16'b01111_010101_01010;
        onion_soup_dim[15][1] = 16'b01111_010101_01010;
        onion_soup_dim[15][2] = 16'b01111_010101_01010;
        onion_soup_dim[15][3] = 16'b01111_010101_01010;
        onion_soup_dim[15][4] = 16'b00110_000111_00000;
        onion_soup_dim[15][5] = 16'b00111_000111_00000;
        onion_soup_dim[15][6] = 16'b01000_001001_00001;
        onion_soup_dim[15][7] = 16'b00110_000111_00000;
        onion_soup_dim[15][8] = 16'b01100_010000_00011;
        onion_soup_dim[15][9] = 16'b01101_010011_00101;
        onion_soup_dim[15][10] = 16'b01100_010001_00011;
        onion_soup_dim[15][11] = 16'b00101_000101_00000;
        onion_soup_dim[15][12] = 16'b00110_000111_00000;
        onion_soup_dim[15][13] = 16'b00101_000110_00000;
        onion_soup_dim[15][14] = 16'b01000_001001_00001;
        onion_soup_dim[15][15] = 16'b00100_000100_00000;
        onion_soup_dim[15][16] = 16'b00111_001000_00001;
        onion_soup_dim[15][17] = 16'b01000_001001_00001;
        onion_soup_dim[15][18] = 16'b00110_000111_00000;
        onion_soup_dim[15][19] = 16'b00111_001000_00000;
        onion_soup_dim[15][20] = 16'b00111_001000_00000;
        onion_soup_dim[15][21] = 16'b00101_000101_00000;
        onion_soup_dim[15][22] = 16'b00111_001000_00001;
        onion_soup_dim[15][23] = 16'b00110_000111_00000;
        onion_soup_dim[15][24] = 16'b00101_000101_00000;
        onion_soup_dim[15][25] = 16'b00111_001000_00000;
        onion_soup_dim[15][26] = 16'b00111_001000_00001;
        onion_soup_dim[15][27] = 16'b01000_001001_00001;
        onion_soup_dim[15][28] = 16'b01111_010101_01010;
        onion_soup_dim[15][29] = 16'b01111_010101_01010;
        onion_soup_dim[15][30] = 16'b01111_010101_01010;
        onion_soup_dim[15][31] = 16'b01111_010101_01010;
        onion_soup_dim[16][0] = 16'b01111_010101_01010;
        onion_soup_dim[16][1] = 16'b01111_010101_01010;
        onion_soup_dim[16][2] = 16'b01111_010101_01010;
        onion_soup_dim[16][3] = 16'b01111_010101_01010;
        onion_soup_dim[16][4] = 16'b01000_001010_00001;
        onion_soup_dim[16][5] = 16'b01001_001100_00001;
        onion_soup_dim[16][6] = 16'b00101_000110_00000;
        onion_soup_dim[16][7] = 16'b00110_000110_00000;
        onion_soup_dim[16][8] = 16'b00111_001000_00000;
        onion_soup_dim[16][9] = 16'b00110_000111_00000;
        onion_soup_dim[16][10] = 16'b00101_000101_00000;
        onion_soup_dim[16][11] = 16'b00111_001000_00000;
        onion_soup_dim[16][12] = 16'b00111_001000_00000;
        onion_soup_dim[16][13] = 16'b00101_000110_00000;
        onion_soup_dim[16][14] = 16'b00110_000111_00001;
        onion_soup_dim[16][15] = 16'b01011_010000_00011;
        onion_soup_dim[16][16] = 16'b01101_010011_00100;
        onion_soup_dim[16][17] = 16'b01000_001001_00001;
        onion_soup_dim[16][18] = 16'b00110_000111_00000;
        onion_soup_dim[16][19] = 16'b00101_000101_00000;
        onion_soup_dim[16][20] = 16'b00101_000100_00000;
        onion_soup_dim[16][21] = 16'b01010_001100_00010;
        onion_soup_dim[16][22] = 16'b01011_010000_00100;
        onion_soup_dim[16][23] = 16'b01101_010110_00111;
        onion_soup_dim[16][24] = 16'b00111_000111_00000;
        onion_soup_dim[16][25] = 16'b00110_000110_00000;
        onion_soup_dim[16][26] = 16'b01000_001010_00001;
        onion_soup_dim[16][27] = 16'b00111_001000_00000;
        onion_soup_dim[16][28] = 16'b01111_010101_01010;
        onion_soup_dim[16][29] = 16'b01111_010101_01010;
        onion_soup_dim[16][30] = 16'b01111_010101_01010;
        onion_soup_dim[16][31] = 16'b01111_010101_01010;
        onion_soup_dim[17][0] = 16'b01111_010101_01010;
        onion_soup_dim[17][1] = 16'b01111_010101_01010;
        onion_soup_dim[17][2] = 16'b01111_010101_01010;
        onion_soup_dim[17][3] = 16'b01111_010101_01010;
        onion_soup_dim[17][4] = 16'b00110_000111_00000;
        onion_soup_dim[17][5] = 16'b01000_001010_00001;
        onion_soup_dim[17][6] = 16'b00101_000101_00000;
        onion_soup_dim[17][7] = 16'b00101_000101_00000;
        onion_soup_dim[17][8] = 16'b00110_000110_00000;
        onion_soup_dim[17][9] = 16'b00111_000111_00000;
        onion_soup_dim[17][10] = 16'b01001_001011_00001;
        onion_soup_dim[17][11] = 16'b01001_001011_00001;
        onion_soup_dim[17][12] = 16'b00111_000111_00000;
        onion_soup_dim[17][13] = 16'b00110_000111_00000;
        onion_soup_dim[17][14] = 16'b01000_001010_00001;
        onion_soup_dim[17][15] = 16'b00111_001000_00001;
        onion_soup_dim[17][16] = 16'b00111_001000_00001;
        onion_soup_dim[17][17] = 16'b01000_001010_00001;
        onion_soup_dim[17][18] = 16'b00110_000110_00000;
        onion_soup_dim[17][19] = 16'b01000_001010_00001;
        onion_soup_dim[17][20] = 16'b00111_001000_00001;
        onion_soup_dim[17][21] = 16'b00110_000111_00000;
        onion_soup_dim[17][22] = 16'b00111_000111_00000;
        onion_soup_dim[17][23] = 16'b00101_000101_00000;
        onion_soup_dim[17][24] = 16'b00101_000110_00000;
        onion_soup_dim[17][25] = 16'b00111_001000_00001;
        onion_soup_dim[17][26] = 16'b00111_001001_00001;
        onion_soup_dim[17][27] = 16'b01000_001011_00001;
        onion_soup_dim[17][28] = 16'b01111_010101_01010;
        onion_soup_dim[17][29] = 16'b01111_010101_01010;
        onion_soup_dim[17][30] = 16'b01111_010101_01010;
        onion_soup_dim[17][31] = 16'b01111_010101_01010;
        onion_soup_dim[18][0] = 16'b01111_010101_01010;
        onion_soup_dim[18][1] = 16'b01111_010101_01010;
        onion_soup_dim[18][2] = 16'b01111_010101_01010;
        onion_soup_dim[18][3] = 16'b01111_010101_01010;
        onion_soup_dim[18][4] = 16'b00111_000111_00001;
        onion_soup_dim[18][5] = 16'b01011_010000_00011;
        onion_soup_dim[18][6] = 16'b00100_000100_00000;
        onion_soup_dim[18][7] = 16'b00101_000110_00000;
        onion_soup_dim[18][8] = 16'b00101_000101_00000;
        onion_soup_dim[18][9] = 16'b00101_000101_00000;
        onion_soup_dim[18][10] = 16'b00111_001000_00001;
        onion_soup_dim[18][11] = 16'b01101_010100_00110;
        onion_soup_dim[18][12] = 16'b01001_001100_00010;
        onion_soup_dim[18][13] = 16'b00110_000110_00000;
        onion_soup_dim[18][14] = 16'b00111_001000_00001;
        onion_soup_dim[18][15] = 16'b01000_001010_00001;
        onion_soup_dim[18][16] = 16'b00111_001000_00000;
        onion_soup_dim[18][17] = 16'b00110_000111_00000;
        onion_soup_dim[18][18] = 16'b01000_001100_00011;
        onion_soup_dim[18][19] = 16'b01011_010000_00011;
        onion_soup_dim[18][20] = 16'b01011_010000_00100;
        onion_soup_dim[18][21] = 16'b00110_000110_00000;
        onion_soup_dim[18][22] = 16'b00110_000110_00000;
        onion_soup_dim[18][23] = 16'b00101_000101_00000;
        onion_soup_dim[18][24] = 16'b00111_000111_00000;
        onion_soup_dim[18][25] = 16'b01000_001010_00001;
        onion_soup_dim[18][26] = 16'b01001_001100_00010;
        onion_soup_dim[18][27] = 16'b01011_010000_00011;
        onion_soup_dim[18][28] = 16'b01111_010101_01010;
        onion_soup_dim[18][29] = 16'b01111_010101_01010;
        onion_soup_dim[18][30] = 16'b01111_010101_01010;
        onion_soup_dim[18][31] = 16'b01111_010101_01010;
        onion_soup_dim[19][0] = 16'b01111_010101_01010;
        onion_soup_dim[19][1] = 16'b01111_010101_01010;
        onion_soup_dim[19][2] = 16'b01111_010101_01010;
        onion_soup_dim[19][3] = 16'b01111_010101_01010;
        onion_soup_dim[19][4] = 16'b01111_010101_01010;
        onion_soup_dim[19][5] = 16'b00110_000111_00001;
        onion_soup_dim[19][6] = 16'b01010_001110_00010;
        onion_soup_dim[19][7] = 16'b00101_000101_00000;
        onion_soup_dim[19][8] = 16'b00110_000111_00000;
        onion_soup_dim[19][9] = 16'b00101_000101_00000;
        onion_soup_dim[19][10] = 16'b00101_000101_00000;
        onion_soup_dim[19][11] = 16'b00111_001000_00001;
        onion_soup_dim[19][12] = 16'b01000_001001_00001;
        onion_soup_dim[19][13] = 16'b00101_000110_00000;
        onion_soup_dim[19][14] = 16'b00101_000101_00000;
        onion_soup_dim[19][15] = 16'b00101_000101_00000;
        onion_soup_dim[19][16] = 16'b00101_000101_00000;
        onion_soup_dim[19][17] = 16'b00111_001000_00000;
        onion_soup_dim[19][18] = 16'b00110_000110_00000;
        onion_soup_dim[19][19] = 16'b00110_000110_00000;
        onion_soup_dim[19][20] = 16'b00101_000101_00000;
        onion_soup_dim[19][21] = 16'b00100_000100_00000;
        onion_soup_dim[19][22] = 16'b00101_000101_00000;
        onion_soup_dim[19][23] = 16'b00101_000101_00000;
        onion_soup_dim[19][24] = 16'b00110_000110_00000;
        onion_soup_dim[19][25] = 16'b01011_001110_00010;
        onion_soup_dim[19][26] = 16'b01001_001100_00010;
        onion_soup_dim[19][27] = 16'b01111_010101_01010;
        onion_soup_dim[19][28] = 16'b01111_010101_01010;
        onion_soup_dim[19][29] = 16'b01111_010101_01010;
        onion_soup_dim[19][30] = 16'b01111_010101_01010;
        onion_soup_dim[19][31] = 16'b01111_010101_01010;
        onion_soup_dim[20][0] = 16'b01111_010101_01010;
        onion_soup_dim[20][1] = 16'b01111_010101_01010;
        onion_soup_dim[20][2] = 16'b01111_010101_01010;
        onion_soup_dim[20][3] = 16'b01111_010101_01010;
        onion_soup_dim[20][4] = 16'b01111_010101_01010;
        onion_soup_dim[20][5] = 16'b01100_010001_00100;
        onion_soup_dim[20][6] = 16'b00110_001000_00001;
        onion_soup_dim[20][7] = 16'b01001_001101_00010;
        onion_soup_dim[20][8] = 16'b00111_001000_00001;
        onion_soup_dim[20][9] = 16'b00111_001001_00001;
        onion_soup_dim[20][10] = 16'b00110_000111_00000;
        onion_soup_dim[20][11] = 16'b01000_001001_00001;
        onion_soup_dim[20][12] = 16'b00110_000111_00000;
        onion_soup_dim[20][13] = 16'b00111_001000_00000;
        onion_soup_dim[20][14] = 16'b00100_000100_00000;
        onion_soup_dim[20][15] = 16'b00101_000110_00000;
        onion_soup_dim[20][16] = 16'b00101_000110_00000;
        onion_soup_dim[20][17] = 16'b00110_000111_00000;
        onion_soup_dim[20][18] = 16'b00110_000111_00000;
        onion_soup_dim[20][19] = 16'b00110_000111_00000;
        onion_soup_dim[20][20] = 16'b00111_000111_00000;
        onion_soup_dim[20][21] = 16'b00111_001000_00001;
        onion_soup_dim[20][22] = 16'b01000_001001_00001;
        onion_soup_dim[20][23] = 16'b00111_001000_00001;
        onion_soup_dim[20][24] = 16'b01001_001100_00010;
        onion_soup_dim[20][25] = 16'b01001_001011_00001;
        onion_soup_dim[20][26] = 16'b01100_010001_00011;
        onion_soup_dim[20][27] = 16'b01111_010101_01010;
        onion_soup_dim[20][28] = 16'b01111_010101_01010;
        onion_soup_dim[20][29] = 16'b01111_010101_01010;
        onion_soup_dim[20][30] = 16'b01111_010101_01010;
        onion_soup_dim[20][31] = 16'b01111_010101_01010;
        onion_soup_dim[21][0] = 16'b01111_010101_01010;
        onion_soup_dim[21][1] = 16'b01111_010101_01010;
        onion_soup_dim[21][2] = 16'b01111_010101_01010;
        onion_soup_dim[21][3] = 16'b01111_010101_01010;
        onion_soup_dim[21][4] = 16'b01111_010101_01010;
        onion_soup_dim[21][5] = 16'b01111_010101_01010;
        onion_soup_dim[21][6] = 16'b01001_001100_00010;
        onion_soup_dim[21][7] = 16'b01000_001010_00001;
        onion_soup_dim[21][8] = 16'b01000_001001_00001;
        onion_soup_dim[21][9] = 16'b01011_001110_00011;
        onion_soup_dim[21][10] = 16'b01000_001010_00001;
        onion_soup_dim[21][11] = 16'b01000_001001_00001;
        onion_soup_dim[21][12] = 16'b01010_001101_00010;
        onion_soup_dim[21][13] = 16'b01000_001010_00001;
        onion_soup_dim[21][14] = 16'b01000_001001_00001;
        onion_soup_dim[21][15] = 16'b01011_001111_00011;
        onion_soup_dim[21][16] = 16'b01010_001101_00010;
        onion_soup_dim[21][17] = 16'b01000_001011_00001;
        onion_soup_dim[21][18] = 16'b01010_001110_00010;
        onion_soup_dim[21][19] = 16'b01001_001011_00010;
        onion_soup_dim[21][20] = 16'b01000_001010_00001;
        onion_soup_dim[21][21] = 16'b01010_001101_00010;
        onion_soup_dim[21][22] = 16'b01011_001110_00011;
        onion_soup_dim[21][23] = 16'b01010_001100_00010;
        onion_soup_dim[21][24] = 16'b01000_001011_00001;
        onion_soup_dim[21][25] = 16'b01010_001110_00011;
        onion_soup_dim[21][26] = 16'b01001_001110_00011;
        onion_soup_dim[21][27] = 16'b01111_010101_01010;
        onion_soup_dim[21][28] = 16'b01111_010101_01010;
        onion_soup_dim[21][29] = 16'b01111_010101_01010;
        onion_soup_dim[21][30] = 16'b01111_010101_01010;
        onion_soup_dim[21][31] = 16'b01111_010101_01010;
        onion_soup_dim[22][0] = 16'b01111_010101_01010;
        onion_soup_dim[22][1] = 16'b01111_010101_01010;
        onion_soup_dim[22][2] = 16'b01111_010101_01010;
        onion_soup_dim[22][3] = 16'b01111_010101_01010;
        onion_soup_dim[22][4] = 16'b01111_010101_01010;
        onion_soup_dim[22][5] = 16'b01111_010101_01010;
        onion_soup_dim[22][6] = 16'b01111_010101_01010;
        onion_soup_dim[22][7] = 16'b01111_010101_01010;
        onion_soup_dim[22][8] = 16'b01001_001100_00010;
        onion_soup_dim[22][9] = 16'b00111_001001_00001;
        onion_soup_dim[22][10] = 16'b01010_001101_00010;
        onion_soup_dim[22][11] = 16'b01010_001100_00010;
        onion_soup_dim[22][12] = 16'b01001_001100_00010;
        onion_soup_dim[22][13] = 16'b01010_001100_00010;
        onion_soup_dim[22][14] = 16'b01100_010001_00100;
        onion_soup_dim[22][15] = 16'b01010_001101_00010;
        onion_soup_dim[22][16] = 16'b01100_010001_00100;
        onion_soup_dim[22][17] = 16'b01101_010011_00101;
        onion_soup_dim[22][18] = 16'b01000_001010_00001;
        onion_soup_dim[22][19] = 16'b01100_010001_00100;
        onion_soup_dim[22][20] = 16'b01011_001111_00011;
        onion_soup_dim[22][21] = 16'b01000_001010_00001;
        onion_soup_dim[22][22] = 16'b01001_001011_00001;
        onion_soup_dim[22][23] = 16'b01011_010000_00011;
        onion_soup_dim[22][24] = 16'b01111_010101_01010;
        onion_soup_dim[22][25] = 16'b01111_010101_01010;
        onion_soup_dim[22][26] = 16'b01111_010101_01010;
        onion_soup_dim[22][27] = 16'b01111_010101_01010;
        onion_soup_dim[22][28] = 16'b01111_010101_01010;
        onion_soup_dim[22][29] = 16'b01111_010101_01010;
        onion_soup_dim[22][30] = 16'b01111_010101_01010;
        onion_soup_dim[22][31] = 16'b01111_010101_01010;
        onion_soup_dim[23][0] = 16'b01111_010101_01010;
        onion_soup_dim[23][1] = 16'b01111_010101_01010;
        onion_soup_dim[23][2] = 16'b01111_010101_01010;
        onion_soup_dim[23][3] = 16'b01111_010101_01010;
        onion_soup_dim[23][4] = 16'b01111_010101_01010;
        onion_soup_dim[23][5] = 16'b01111_010101_01010;
        onion_soup_dim[23][6] = 16'b01111_010101_01010;
        onion_soup_dim[23][7] = 16'b01111_010101_01010;
        onion_soup_dim[23][8] = 16'b01111_010101_01010;
        onion_soup_dim[23][9] = 16'b01111_010101_01010;
        onion_soup_dim[23][10] = 16'b01101_010101_00110;
        onion_soup_dim[23][11] = 16'b01100_010010_00101;
        onion_soup_dim[23][12] = 16'b00111_001000_00001;
        onion_soup_dim[23][13] = 16'b01001_001011_00001;
        onion_soup_dim[23][14] = 16'b01001_001100_00010;
        onion_soup_dim[23][15] = 16'b01010_001110_00010;
        onion_soup_dim[23][16] = 16'b01001_001011_00010;
        onion_soup_dim[23][17] = 16'b01001_001100_00010;
        onion_soup_dim[23][18] = 16'b01100_010001_00011;
        onion_soup_dim[23][19] = 16'b01010_001101_00010;
        onion_soup_dim[23][20] = 16'b01001_001011_00010;
        onion_soup_dim[23][21] = 16'b01101_010101_00111;
        onion_soup_dim[23][22] = 16'b01100_010010_00101;
        onion_soup_dim[23][23] = 16'b01111_010101_01010;
        onion_soup_dim[23][24] = 16'b01111_010101_01010;
        onion_soup_dim[23][25] = 16'b01111_010101_01010;
        onion_soup_dim[23][26] = 16'b01111_010101_01010;
        onion_soup_dim[23][27] = 16'b01111_010101_01010;
        onion_soup_dim[23][28] = 16'b01111_010101_01010;
        onion_soup_dim[23][29] = 16'b01111_010101_01010;
        onion_soup_dim[23][30] = 16'b01111_010101_01010;
        onion_soup_dim[23][31] = 16'b01111_010101_01010;
        onion_soup_dim[24][0] = 16'b01111_010101_01010;
        onion_soup_dim[24][1] = 16'b01111_010101_01010;
        onion_soup_dim[24][2] = 16'b01111_010101_01010;
        onion_soup_dim[24][3] = 16'b01111_010101_01010;
        onion_soup_dim[24][4] = 16'b01111_010101_01010;
        onion_soup_dim[24][5] = 16'b01111_010101_01010;
        onion_soup_dim[24][6] = 16'b01111_010101_01010;
        onion_soup_dim[24][7] = 16'b01111_010101_01010;
        onion_soup_dim[24][8] = 16'b01111_010101_01010;
        onion_soup_dim[24][9] = 16'b01111_010101_01010;
        onion_soup_dim[24][10] = 16'b01111_010101_01010;
        onion_soup_dim[24][11] = 16'b01111_010101_01010;
        onion_soup_dim[24][12] = 16'b01111_010101_01010;
        onion_soup_dim[24][13] = 16'b01111_010101_01010;
        onion_soup_dim[24][14] = 16'b01111_010101_01010;
        onion_soup_dim[24][15] = 16'b01111_010101_01010;
        onion_soup_dim[24][16] = 16'b01111_010101_01010;
        onion_soup_dim[24][17] = 16'b01111_010101_01010;
        onion_soup_dim[24][18] = 16'b01111_010101_01010;
        onion_soup_dim[24][19] = 16'b01111_010101_01010;
        onion_soup_dim[24][20] = 16'b01111_010101_01010;
        onion_soup_dim[24][21] = 16'b01111_010101_01010;
        onion_soup_dim[24][22] = 16'b01111_010101_01010;
        onion_soup_dim[24][23] = 16'b01111_010101_01010;
        onion_soup_dim[24][24] = 16'b01111_010101_01010;
        onion_soup_dim[24][25] = 16'b01111_010101_01010;
        onion_soup_dim[24][26] = 16'b01111_010101_01010;
        onion_soup_dim[24][27] = 16'b01111_010101_01010;
        onion_soup_dim[24][28] = 16'b01111_010101_01010;
        onion_soup_dim[24][29] = 16'b01111_010101_01010;
        onion_soup_dim[24][30] = 16'b01111_010101_01010;
        onion_soup_dim[24][31] = 16'b01111_010101_01010;
        onion_soup_dim[25][0] = 16'b01111_010101_01010;
        onion_soup_dim[25][1] = 16'b01111_010101_01010;
        onion_soup_dim[25][2] = 16'b01111_010101_01010;
        onion_soup_dim[25][3] = 16'b01111_010101_01010;
        onion_soup_dim[25][4] = 16'b01111_010101_01010;
        onion_soup_dim[25][5] = 16'b01111_010101_01010;
        onion_soup_dim[25][6] = 16'b01111_010101_01010;
        onion_soup_dim[25][7] = 16'b01111_010101_01010;
        onion_soup_dim[25][8] = 16'b01111_010101_01010;
        onion_soup_dim[25][9] = 16'b01111_010101_01010;
        onion_soup_dim[25][10] = 16'b01111_010101_01010;
        onion_soup_dim[25][11] = 16'b01111_010101_01010;
        onion_soup_dim[25][12] = 16'b01111_010101_01010;
        onion_soup_dim[25][13] = 16'b01111_010101_01010;
        onion_soup_dim[25][14] = 16'b01111_010101_01010;
        onion_soup_dim[25][15] = 16'b01111_010101_01010;
        onion_soup_dim[25][16] = 16'b01111_010101_01010;
        onion_soup_dim[25][17] = 16'b01111_010101_01010;
        onion_soup_dim[25][18] = 16'b01111_010101_01010;
        onion_soup_dim[25][19] = 16'b01111_010101_01010;
        onion_soup_dim[25][20] = 16'b01111_010101_01010;
        onion_soup_dim[25][21] = 16'b01111_010101_01010;
        onion_soup_dim[25][22] = 16'b01111_010101_01010;
        onion_soup_dim[25][23] = 16'b01111_010101_01010;
        onion_soup_dim[25][24] = 16'b01111_010101_01010;
        onion_soup_dim[25][25] = 16'b01111_010101_01010;
        onion_soup_dim[25][26] = 16'b01111_010101_01010;
        onion_soup_dim[25][27] = 16'b01111_010101_01010;
        onion_soup_dim[25][28] = 16'b01111_010101_01010;
        onion_soup_dim[25][29] = 16'b01111_010101_01010;
        onion_soup_dim[25][30] = 16'b01111_010101_01010;
        onion_soup_dim[25][31] = 16'b01111_010101_01010;
        onion_soup_dim[26][0] = 16'b01111_010101_01010;
        onion_soup_dim[26][1] = 16'b01111_010101_01010;
        onion_soup_dim[26][2] = 16'b01111_010101_01010;
        onion_soup_dim[26][3] = 16'b01111_010101_01010;
        onion_soup_dim[26][4] = 16'b01111_010101_01010;
        onion_soup_dim[26][5] = 16'b01111_010101_01010;
        onion_soup_dim[26][6] = 16'b01111_010101_01010;
        onion_soup_dim[26][7] = 16'b01111_010101_01010;
        onion_soup_dim[26][8] = 16'b01111_010101_01010;
        onion_soup_dim[26][9] = 16'b01111_010101_01010;
        onion_soup_dim[26][10] = 16'b01111_010101_01010;
        onion_soup_dim[26][11] = 16'b01111_010101_01010;
        onion_soup_dim[26][12] = 16'b01111_010101_01010;
        onion_soup_dim[26][13] = 16'b01111_010101_01010;
        onion_soup_dim[26][14] = 16'b01111_010101_01010;
        onion_soup_dim[26][15] = 16'b01111_010101_01010;
        onion_soup_dim[26][16] = 16'b01111_010101_01010;
        onion_soup_dim[26][17] = 16'b01111_010101_01010;
        onion_soup_dim[26][18] = 16'b01111_010101_01010;
        onion_soup_dim[26][19] = 16'b01111_010101_01010;
        onion_soup_dim[26][20] = 16'b01111_010101_01010;
        onion_soup_dim[26][21] = 16'b01111_010101_01010;
        onion_soup_dim[26][22] = 16'b01111_010101_01010;
        onion_soup_dim[26][23] = 16'b01111_010101_01010;
        onion_soup_dim[26][24] = 16'b01111_010101_01010;
        onion_soup_dim[26][25] = 16'b01111_010101_01010;
        onion_soup_dim[26][26] = 16'b01111_010101_01010;
        onion_soup_dim[26][27] = 16'b01111_010101_01010;
        onion_soup_dim[26][28] = 16'b01111_010101_01010;
        onion_soup_dim[26][29] = 16'b01111_010101_01010;
        onion_soup_dim[26][30] = 16'b01111_010101_01010;
        onion_soup_dim[26][31] = 16'b01111_010101_01010;
        onion_soup_dim[27][0] = 16'b01111_010101_01010;
        onion_soup_dim[27][1] = 16'b01111_010101_01010;
        onion_soup_dim[27][2] = 16'b01111_010101_01010;
        onion_soup_dim[27][3] = 16'b01111_010101_01010;
        onion_soup_dim[27][4] = 16'b01111_010101_01010;
        onion_soup_dim[27][5] = 16'b01111_010101_01010;
        onion_soup_dim[27][6] = 16'b01111_010101_01010;
        onion_soup_dim[27][7] = 16'b01111_010101_01010;
        onion_soup_dim[27][8] = 16'b01111_010101_01010;
        onion_soup_dim[27][9] = 16'b01111_010101_01010;
        onion_soup_dim[27][10] = 16'b01111_010101_01010;
        onion_soup_dim[27][11] = 16'b01111_010101_01010;
        onion_soup_dim[27][12] = 16'b01111_010101_01010;
        onion_soup_dim[27][13] = 16'b01111_010101_01010;
        onion_soup_dim[27][14] = 16'b01111_010101_01010;
        onion_soup_dim[27][15] = 16'b01111_010101_01010;
        onion_soup_dim[27][16] = 16'b01111_010101_01010;
        onion_soup_dim[27][17] = 16'b01111_010101_01010;
        onion_soup_dim[27][18] = 16'b01111_010101_01010;
        onion_soup_dim[27][19] = 16'b01111_010101_01010;
        onion_soup_dim[27][20] = 16'b01111_010101_01010;
        onion_soup_dim[27][21] = 16'b01111_010101_01010;
        onion_soup_dim[27][22] = 16'b01111_010101_01010;
        onion_soup_dim[27][23] = 16'b01111_010101_01010;
        onion_soup_dim[27][24] = 16'b01111_010101_01010;
        onion_soup_dim[27][25] = 16'b01111_010101_01010;
        onion_soup_dim[27][26] = 16'b01111_010101_01010;
        onion_soup_dim[27][27] = 16'b01111_010101_01010;
        onion_soup_dim[27][28] = 16'b01111_010101_01010;
        onion_soup_dim[27][29] = 16'b01111_010101_01010;
        onion_soup_dim[27][30] = 16'b01111_010101_01010;
        onion_soup_dim[27][31] = 16'b01111_010101_01010;
        onion_soup_dim[28][0] = 16'b01111_010101_01010;
        onion_soup_dim[28][1] = 16'b01111_010101_01010;
        onion_soup_dim[28][2] = 16'b01111_010101_01010;
        onion_soup_dim[28][3] = 16'b01111_010101_01010;
        onion_soup_dim[28][4] = 16'b01111_010101_01010;
        onion_soup_dim[28][5] = 16'b01111_010101_01010;
        onion_soup_dim[28][6] = 16'b01111_010101_01010;
        onion_soup_dim[28][7] = 16'b01111_010101_01010;
        onion_soup_dim[28][8] = 16'b01111_010101_01010;
        onion_soup_dim[28][9] = 16'b01111_010101_01010;
        onion_soup_dim[28][10] = 16'b01111_010101_01010;
        onion_soup_dim[28][11] = 16'b01111_010101_01010;
        onion_soup_dim[28][12] = 16'b01111_010101_01010;
        onion_soup_dim[28][13] = 16'b01111_010101_01010;
        onion_soup_dim[28][14] = 16'b01111_010101_01010;
        onion_soup_dim[28][15] = 16'b01111_010101_01010;
        onion_soup_dim[28][16] = 16'b01111_010101_01010;
        onion_soup_dim[28][17] = 16'b01111_010101_01010;
        onion_soup_dim[28][18] = 16'b01111_010101_01010;
        onion_soup_dim[28][19] = 16'b01111_010101_01010;
        onion_soup_dim[28][20] = 16'b01111_010101_01010;
        onion_soup_dim[28][21] = 16'b01111_010101_01010;
        onion_soup_dim[28][22] = 16'b01111_010101_01010;
        onion_soup_dim[28][23] = 16'b01111_010101_01010;
        onion_soup_dim[28][24] = 16'b01111_010101_01010;
        onion_soup_dim[28][25] = 16'b01111_010101_01010;
        onion_soup_dim[28][26] = 16'b01111_010101_01010;
        onion_soup_dim[28][27] = 16'b01111_010101_01010;
        onion_soup_dim[28][28] = 16'b01111_010101_01010;
        onion_soup_dim[28][29] = 16'b01111_010101_01010;
        onion_soup_dim[28][30] = 16'b01111_010101_01010;
        onion_soup_dim[28][31] = 16'b01111_010101_01010;
        onion_soup_dim[29][0] = 16'b01111_010101_01010;
        onion_soup_dim[29][1] = 16'b01111_010101_01010;
        onion_soup_dim[29][2] = 16'b01111_010101_01010;
        onion_soup_dim[29][3] = 16'b01111_010101_01010;
        onion_soup_dim[29][4] = 16'b01111_010101_01010;
        onion_soup_dim[29][5] = 16'b01111_010101_01010;
        onion_soup_dim[29][6] = 16'b01111_010101_01010;
        onion_soup_dim[29][7] = 16'b01111_010101_01010;
        onion_soup_dim[29][8] = 16'b01111_010101_01010;
        onion_soup_dim[29][9] = 16'b01111_010101_01010;
        onion_soup_dim[29][10] = 16'b01111_010101_01010;
        onion_soup_dim[29][11] = 16'b01111_010101_01010;
        onion_soup_dim[29][12] = 16'b01111_010101_01010;
        onion_soup_dim[29][13] = 16'b01111_010101_01010;
        onion_soup_dim[29][14] = 16'b01111_010101_01010;
        onion_soup_dim[29][15] = 16'b01111_010101_01010;
        onion_soup_dim[29][16] = 16'b01111_010101_01010;
        onion_soup_dim[29][17] = 16'b01111_010101_01010;
        onion_soup_dim[29][18] = 16'b01111_010101_01010;
        onion_soup_dim[29][19] = 16'b01111_010101_01010;
        onion_soup_dim[29][20] = 16'b01111_010101_01010;
        onion_soup_dim[29][21] = 16'b01111_010101_01010;
        onion_soup_dim[29][22] = 16'b01111_010101_01010;
        onion_soup_dim[29][23] = 16'b01111_010101_01010;
        onion_soup_dim[29][24] = 16'b01111_010101_01010;
        onion_soup_dim[29][25] = 16'b01111_010101_01010;
        onion_soup_dim[29][26] = 16'b01111_010101_01010;
        onion_soup_dim[29][27] = 16'b01111_010101_01010;
        onion_soup_dim[29][28] = 16'b01111_010101_01010;
        onion_soup_dim[29][29] = 16'b01111_010101_01010;
        onion_soup_dim[29][30] = 16'b01111_010101_01010;
        onion_soup_dim[29][31] = 16'b01111_010101_01010;
        onion_soup_dim[30][0] = 16'b01111_010101_01010;
        onion_soup_dim[30][1] = 16'b01111_010101_01010;
        onion_soup_dim[30][2] = 16'b01111_010101_01010;
        onion_soup_dim[30][3] = 16'b01111_010101_01010;
        onion_soup_dim[30][4] = 16'b01111_010101_01010;
        onion_soup_dim[30][5] = 16'b01111_010101_01010;
        onion_soup_dim[30][6] = 16'b01111_010101_01010;
        onion_soup_dim[30][7] = 16'b01111_010101_01010;
        onion_soup_dim[30][8] = 16'b01111_010101_01010;
        onion_soup_dim[30][9] = 16'b01111_010101_01010;
        onion_soup_dim[30][10] = 16'b01111_010101_01010;
        onion_soup_dim[30][11] = 16'b01111_010101_01010;
        onion_soup_dim[30][12] = 16'b01111_010101_01010;
        onion_soup_dim[30][13] = 16'b01111_010101_01010;
        onion_soup_dim[30][14] = 16'b01111_010101_01010;
        onion_soup_dim[30][15] = 16'b01111_010101_01010;
        onion_soup_dim[30][16] = 16'b01111_010101_01010;
        onion_soup_dim[30][17] = 16'b01111_010101_01010;
        onion_soup_dim[30][18] = 16'b01111_010101_01010;
        onion_soup_dim[30][19] = 16'b01111_010101_01010;
        onion_soup_dim[30][20] = 16'b01111_010101_01010;
        onion_soup_dim[30][21] = 16'b01111_010101_01010;
        onion_soup_dim[30][22] = 16'b01111_010101_01010;
        onion_soup_dim[30][23] = 16'b01111_010101_01010;
        onion_soup_dim[30][24] = 16'b01111_010101_01010;
        onion_soup_dim[30][25] = 16'b01111_010101_01010;
        onion_soup_dim[30][26] = 16'b01111_010101_01010;
        onion_soup_dim[30][27] = 16'b01111_010101_01010;
        onion_soup_dim[30][28] = 16'b01111_010101_01010;
        onion_soup_dim[30][29] = 16'b01111_010101_01010;
        onion_soup_dim[30][30] = 16'b01111_010101_01010;
        onion_soup_dim[30][31] = 16'b01111_010101_01010;
        onion_soup_dim[31][0] = 16'b01111_010101_01010;
        onion_soup_dim[31][1] = 16'b01111_010101_01010;
        onion_soup_dim[31][2] = 16'b01111_010101_01010;
        onion_soup_dim[31][3] = 16'b01111_010101_01010;
        onion_soup_dim[31][4] = 16'b01111_010101_01010;
        onion_soup_dim[31][5] = 16'b01111_010101_01010;
        onion_soup_dim[31][6] = 16'b01111_010101_01010;
        onion_soup_dim[31][7] = 16'b01111_010101_01010;
        onion_soup_dim[31][8] = 16'b01111_010101_01010;
        onion_soup_dim[31][9] = 16'b01111_010101_01010;
        onion_soup_dim[31][10] = 16'b01111_010101_01010;
        onion_soup_dim[31][11] = 16'b01111_010101_01010;
        onion_soup_dim[31][12] = 16'b01111_010101_01010;
        onion_soup_dim[31][13] = 16'b01111_010101_01010;
        onion_soup_dim[31][14] = 16'b01111_010101_01010;
        onion_soup_dim[31][15] = 16'b01111_010101_01010;
        onion_soup_dim[31][16] = 16'b01111_010101_01010;
        onion_soup_dim[31][17] = 16'b01111_010101_01010;
        onion_soup_dim[31][18] = 16'b01111_010101_01010;
        onion_soup_dim[31][19] = 16'b01111_010101_01010;
        onion_soup_dim[31][20] = 16'b01111_010101_01010;
        onion_soup_dim[31][21] = 16'b01111_010101_01010;
        onion_soup_dim[31][22] = 16'b01111_010101_01010;
        onion_soup_dim[31][23] = 16'b01111_010101_01010;
        onion_soup_dim[31][24] = 16'b01111_010101_01010;
        onion_soup_dim[31][25] = 16'b01111_010101_01010;
        onion_soup_dim[31][26] = 16'b01111_010101_01010;
        onion_soup_dim[31][27] = 16'b01111_010101_01010;
        onion_soup_dim[31][28] = 16'b01111_010101_01010;
        onion_soup_dim[31][29] = 16'b01111_010101_01010;
        onion_soup_dim[31][30] = 16'b01111_010101_01010;
        onion_soup_dim[31][31] = 16'b01111_010101_01010;
        
        
        
                
        tomato_soup_dim[0][0] = 16'b01011_011111_01010;
        tomato_soup_dim[0][1] = 16'b01011_011111_01010;
        tomato_soup_dim[0][2] = 16'b01011_011111_01010;
        tomato_soup_dim[0][3] = 16'b01011_011111_01010;
        tomato_soup_dim[0][4] = 16'b01011_011111_01010;
        tomato_soup_dim[0][5] = 16'b01011_011111_01010;
        tomato_soup_dim[0][6] = 16'b01011_011111_01010;
        tomato_soup_dim[0][7] = 16'b01011_011111_01010;
        tomato_soup_dim[0][8] = 16'b01011_011111_01010;
        tomato_soup_dim[0][9] = 16'b01011_011111_01010;
        tomato_soup_dim[0][10] = 16'b01011_011111_01010;
        tomato_soup_dim[0][11] = 16'b01011_011111_01010;
        tomato_soup_dim[0][12] = 16'b01011_011111_01010;
        tomato_soup_dim[0][13] = 16'b01011_011111_01010;
        tomato_soup_dim[0][14] = 16'b01011_011111_01010;
        tomato_soup_dim[0][15] = 16'b01011_011111_01010;
        tomato_soup_dim[0][16] = 16'b01011_011111_01010;
        tomato_soup_dim[0][17] = 16'b01011_011111_01010;
        tomato_soup_dim[0][18] = 16'b01011_011111_01010;
        tomato_soup_dim[0][19] = 16'b01011_011111_01010;
        tomato_soup_dim[0][20] = 16'b01011_011111_01010;
        tomato_soup_dim[0][21] = 16'b01011_011111_01010;
        tomato_soup_dim[0][22] = 16'b01011_011111_01010;
        tomato_soup_dim[0][23] = 16'b01011_011111_01010;
        tomato_soup_dim[0][24] = 16'b01011_011111_01010;
        tomato_soup_dim[0][25] = 16'b01011_011111_01010;
        tomato_soup_dim[0][26] = 16'b01011_011111_01010;
        tomato_soup_dim[0][27] = 16'b01011_011111_01010;
        tomato_soup_dim[0][28] = 16'b01011_011111_01010;
        tomato_soup_dim[0][29] = 16'b01011_011111_01010;
        tomato_soup_dim[0][30] = 16'b01011_011111_01010;
        tomato_soup_dim[0][31] = 16'b01011_011111_01010;
        tomato_soup_dim[1][0] = 16'b01011_011111_01010;
        tomato_soup_dim[1][1] = 16'b01011_011111_01010;
        tomato_soup_dim[1][2] = 16'b01011_011111_01010;
        tomato_soup_dim[1][3] = 16'b01011_011111_01010;
        tomato_soup_dim[1][4] = 16'b01011_011111_01010;
        tomato_soup_dim[1][5] = 16'b01011_011111_01010;
        tomato_soup_dim[1][6] = 16'b01011_011111_01010;
        tomato_soup_dim[1][7] = 16'b01011_011111_01010;
        tomato_soup_dim[1][8] = 16'b01011_011111_01010;
        tomato_soup_dim[1][9] = 16'b01011_011111_01010;
        tomato_soup_dim[1][10] = 16'b01011_011111_01010;
        tomato_soup_dim[1][11] = 16'b01011_011111_01010;
        tomato_soup_dim[1][12] = 16'b01011_011111_01010;
        tomato_soup_dim[1][13] = 16'b01011_011111_01010;
        tomato_soup_dim[1][14] = 16'b01011_011111_01010;
        tomato_soup_dim[1][15] = 16'b01011_011111_01010;
        tomato_soup_dim[1][16] = 16'b01011_011111_01010;
        tomato_soup_dim[1][17] = 16'b01011_011111_01010;
        tomato_soup_dim[1][18] = 16'b01011_011111_01010;
        tomato_soup_dim[1][19] = 16'b01011_011111_01010;
        tomato_soup_dim[1][20] = 16'b01011_011111_01010;
        tomato_soup_dim[1][21] = 16'b01011_011111_01010;
        tomato_soup_dim[1][22] = 16'b01011_011111_01010;
        tomato_soup_dim[1][23] = 16'b01011_011111_01010;
        tomato_soup_dim[1][24] = 16'b01011_011111_01010;
        tomato_soup_dim[1][25] = 16'b01011_011111_01010;
        tomato_soup_dim[1][26] = 16'b01011_011111_01010;
        tomato_soup_dim[1][27] = 16'b01011_011111_01010;
        tomato_soup_dim[1][28] = 16'b01011_011111_01010;
        tomato_soup_dim[1][29] = 16'b01011_011111_01010;
        tomato_soup_dim[1][30] = 16'b01011_011111_01010;
        tomato_soup_dim[1][31] = 16'b01011_011111_01010;
        tomato_soup_dim[2][0] = 16'b01011_011111_01010;
        tomato_soup_dim[2][1] = 16'b01011_011111_01010;
        tomato_soup_dim[2][2] = 16'b01011_011111_01010;
        tomato_soup_dim[2][3] = 16'b01011_011111_01010;
        tomato_soup_dim[2][4] = 16'b01011_011111_01010;
        tomato_soup_dim[2][5] = 16'b01011_011111_01010;
        tomato_soup_dim[2][6] = 16'b01011_011111_01010;
        tomato_soup_dim[2][7] = 16'b01011_011111_01010;
        tomato_soup_dim[2][8] = 16'b01011_011111_01010;
        tomato_soup_dim[2][9] = 16'b01011_011111_01010;
        tomato_soup_dim[2][10] = 16'b01011_011111_01010;
        tomato_soup_dim[2][11] = 16'b01011_011111_01010;
        tomato_soup_dim[2][12] = 16'b01011_011111_01010;
        tomato_soup_dim[2][13] = 16'b01011_011111_01010;
        tomato_soup_dim[2][14] = 16'b01011_011111_01010;
        tomato_soup_dim[2][15] = 16'b01011_011111_01010;
        tomato_soup_dim[2][16] = 16'b01011_011111_01010;
        tomato_soup_dim[2][17] = 16'b01011_011111_01010;
        tomato_soup_dim[2][18] = 16'b01011_011111_01010;
        tomato_soup_dim[2][19] = 16'b01011_011111_01010;
        tomato_soup_dim[2][20] = 16'b01011_011111_01010;
        tomato_soup_dim[2][21] = 16'b01011_011111_01010;
        tomato_soup_dim[2][22] = 16'b01011_011111_01010;
        tomato_soup_dim[2][23] = 16'b01011_011111_01010;
        tomato_soup_dim[2][24] = 16'b01011_011111_01010;
        tomato_soup_dim[2][25] = 16'b01011_011111_01010;
        tomato_soup_dim[2][26] = 16'b01011_011111_01010;
        tomato_soup_dim[2][27] = 16'b01011_011111_01010;
        tomato_soup_dim[2][28] = 16'b01011_011111_01010;
        tomato_soup_dim[2][29] = 16'b01011_011111_01010;
        tomato_soup_dim[2][30] = 16'b01011_011111_01010;
        tomato_soup_dim[2][31] = 16'b01011_011111_01010;
        tomato_soup_dim[3][0] = 16'b01011_011111_01010;
        tomato_soup_dim[3][1] = 16'b01011_011111_01010;
        tomato_soup_dim[3][2] = 16'b01011_011111_01010;
        tomato_soup_dim[3][3] = 16'b01011_011111_01010;
        tomato_soup_dim[3][4] = 16'b01011_011111_01010;
        tomato_soup_dim[3][5] = 16'b01011_011111_01010;
        tomato_soup_dim[3][6] = 16'b01011_011111_01010;
        tomato_soup_dim[3][7] = 16'b01011_011111_01010;
        tomato_soup_dim[3][8] = 16'b01011_011111_01010;
        tomato_soup_dim[3][9] = 16'b01011_011111_01010;
        tomato_soup_dim[3][10] = 16'b01011_011111_01010;
        tomato_soup_dim[3][11] = 16'b01011_011111_01010;
        tomato_soup_dim[3][12] = 16'b01011_011111_01010;
        tomato_soup_dim[3][13] = 16'b01011_011111_01010;
        tomato_soup_dim[3][14] = 16'b01011_011111_01010;
        tomato_soup_dim[3][15] = 16'b01011_011111_01010;
        tomato_soup_dim[3][16] = 16'b01011_011111_01010;
        tomato_soup_dim[3][17] = 16'b01011_011111_01010;
        tomato_soup_dim[3][18] = 16'b01011_011111_01010;
        tomato_soup_dim[3][19] = 16'b01011_011111_01010;
        tomato_soup_dim[3][20] = 16'b01011_011111_01010;
        tomato_soup_dim[3][21] = 16'b01011_011111_01010;
        tomato_soup_dim[3][22] = 16'b01011_011111_01010;
        tomato_soup_dim[3][23] = 16'b01011_011111_01010;
        tomato_soup_dim[3][24] = 16'b01011_011111_01010;
        tomato_soup_dim[3][25] = 16'b01011_011111_01010;
        tomato_soup_dim[3][26] = 16'b01011_011111_01010;
        tomato_soup_dim[3][27] = 16'b01011_011111_01010;
        tomato_soup_dim[3][28] = 16'b01011_011111_01010;
        tomato_soup_dim[3][29] = 16'b01011_011111_01010;
        tomato_soup_dim[3][30] = 16'b01011_011111_01010;
        tomato_soup_dim[3][31] = 16'b01011_011111_01010;
        tomato_soup_dim[4][0] = 16'b01011_011111_01010;
        tomato_soup_dim[4][1] = 16'b01011_011111_01010;
        tomato_soup_dim[4][2] = 16'b01011_011111_01010;
        tomato_soup_dim[4][3] = 16'b01011_011111_01010;
        tomato_soup_dim[4][4] = 16'b01011_011111_01010;
        tomato_soup_dim[4][5] = 16'b01011_011111_01010;
        tomato_soup_dim[4][6] = 16'b01011_011111_01010;
        tomato_soup_dim[4][7] = 16'b01011_011111_01010;
        tomato_soup_dim[4][8] = 16'b01011_011111_01010;
        tomato_soup_dim[4][9] = 16'b01011_011111_01010;
        tomato_soup_dim[4][10] = 16'b01011_011111_01010;
        tomato_soup_dim[4][11] = 16'b01100_010100_00110;
        tomato_soup_dim[4][12] = 16'b01100_010100_00110;
        tomato_soup_dim[4][13] = 16'b01100_010011_00110;
        tomato_soup_dim[4][14] = 16'b01100_010100_00110;
        tomato_soup_dim[4][15] = 16'b01100_010100_00110;
        tomato_soup_dim[4][16] = 16'b01100_010100_00110;
        tomato_soup_dim[4][17] = 16'b01100_010100_00110;
        tomato_soup_dim[4][18] = 16'b01100_010100_00110;
        tomato_soup_dim[4][19] = 16'b01100_010100_00110;
        tomato_soup_dim[4][20] = 16'b01011_011111_01010;
        tomato_soup_dim[4][21] = 16'b01011_011111_01010;
        tomato_soup_dim[4][22] = 16'b01011_011111_01010;
        tomato_soup_dim[4][23] = 16'b01011_011111_01010;
        tomato_soup_dim[4][24] = 16'b01011_011111_01010;
        tomato_soup_dim[4][25] = 16'b01011_011111_01010;
        tomato_soup_dim[4][26] = 16'b01011_011111_01010;
        tomato_soup_dim[4][27] = 16'b01011_011111_01010;
        tomato_soup_dim[4][28] = 16'b01011_011111_01010;
        tomato_soup_dim[4][29] = 16'b01011_011111_01010;
        tomato_soup_dim[4][30] = 16'b01011_011111_01010;
        tomato_soup_dim[4][31] = 16'b01011_011111_01010;
        tomato_soup_dim[5][0] = 16'b01011_011111_01010;
        tomato_soup_dim[5][1] = 16'b01011_011111_01010;
        tomato_soup_dim[5][2] = 16'b01011_011111_01010;
        tomato_soup_dim[5][3] = 16'b01011_011111_01010;
        tomato_soup_dim[5][4] = 16'b01011_011111_01010;
        tomato_soup_dim[5][5] = 16'b01011_011111_01010;
        tomato_soup_dim[5][6] = 16'b01011_011111_01010;
        tomato_soup_dim[5][7] = 16'b01011_011111_01010;
        tomato_soup_dim[5][8] = 16'b01011_011111_01010;
        tomato_soup_dim[5][9] = 16'b01100_010100_00110;
        tomato_soup_dim[5][10] = 16'b01100_010100_00110;
        tomato_soup_dim[5][11] = 16'b01100_010100_00110;
        tomato_soup_dim[5][12] = 16'b01100_010101_00111;
        tomato_soup_dim[5][13] = 16'b01100_010101_00110;
        tomato_soup_dim[5][14] = 16'b01100_010101_00111;
        tomato_soup_dim[5][15] = 16'b01101_010110_00111;
        tomato_soup_dim[5][16] = 16'b01100_010101_00111;
        tomato_soup_dim[5][17] = 16'b01101_010101_00111;
        tomato_soup_dim[5][18] = 16'b01101_010101_00111;
        tomato_soup_dim[5][19] = 16'b01100_010101_00111;
        tomato_soup_dim[5][20] = 16'b01100_010100_00110;
        tomato_soup_dim[5][21] = 16'b01100_010100_00110;
        tomato_soup_dim[5][22] = 16'b01011_011111_01010;
        tomato_soup_dim[5][23] = 16'b01011_011111_01010;
        tomato_soup_dim[5][24] = 16'b01011_011111_01010;
        tomato_soup_dim[5][25] = 16'b01011_011111_01010;
        tomato_soup_dim[5][26] = 16'b01011_011111_01010;
        tomato_soup_dim[5][27] = 16'b01011_011111_01010;
        tomato_soup_dim[5][28] = 16'b01011_011111_01010;
        tomato_soup_dim[5][29] = 16'b01011_011111_01010;
        tomato_soup_dim[5][30] = 16'b01011_011111_01010;
        tomato_soup_dim[5][31] = 16'b01011_011111_01010;
        tomato_soup_dim[6][0] = 16'b01011_011111_01010;
        tomato_soup_dim[6][1] = 16'b01011_011111_01010;
        tomato_soup_dim[6][2] = 16'b01011_011111_01010;
        tomato_soup_dim[6][3] = 16'b01011_011111_01010;
        tomato_soup_dim[6][4] = 16'b01011_011111_01010;
        tomato_soup_dim[6][5] = 16'b01011_011111_01010;
        tomato_soup_dim[6][6] = 16'b01011_011111_01010;
        tomato_soup_dim[6][7] = 16'b01100_010100_00110;
        tomato_soup_dim[6][8] = 16'b01100_010100_00110;
        tomato_soup_dim[6][9] = 16'b01100_010101_00111;
        tomato_soup_dim[6][10] = 16'b01101_010101_00111;
        tomato_soup_dim[6][11] = 16'b01101_010101_00111;
        tomato_soup_dim[6][12] = 16'b01101_010101_00111;
        tomato_soup_dim[6][13] = 16'b01100_010101_00111;
        tomato_soup_dim[6][14] = 16'b01100_010101_00111;
        tomato_soup_dim[6][15] = 16'b01100_010101_00110;
        tomato_soup_dim[6][16] = 16'b01100_010101_00110;
        tomato_soup_dim[6][17] = 16'b01100_010100_00110;
        tomato_soup_dim[6][18] = 16'b01100_010101_00111;
        tomato_soup_dim[6][19] = 16'b01100_010101_00111;
        tomato_soup_dim[6][20] = 16'b01101_010101_00111;
        tomato_soup_dim[6][21] = 16'b01100_010101_00110;
        tomato_soup_dim[6][22] = 16'b01100_010100_00110;
        tomato_soup_dim[6][23] = 16'b01100_010100_00110;
        tomato_soup_dim[6][24] = 16'b01011_011111_01010;
        tomato_soup_dim[6][25] = 16'b01011_011111_01010;
        tomato_soup_dim[6][26] = 16'b01011_011111_01010;
        tomato_soup_dim[6][27] = 16'b01011_011111_01010;
        tomato_soup_dim[6][28] = 16'b01011_011111_01010;
        tomato_soup_dim[6][29] = 16'b01011_011111_01010;
        tomato_soup_dim[6][30] = 16'b01011_011111_01010;
        tomato_soup_dim[6][31] = 16'b01011_011111_01010;
        tomato_soup_dim[7][0] = 16'b01011_011111_01010;
        tomato_soup_dim[7][1] = 16'b01011_011111_01010;
        tomato_soup_dim[7][2] = 16'b01011_011111_01010;
        tomato_soup_dim[7][3] = 16'b01011_011111_01010;
        tomato_soup_dim[7][4] = 16'b01011_011111_01010;
        tomato_soup_dim[7][5] = 16'b01011_011111_01010;
        tomato_soup_dim[7][6] = 16'b01100_010100_00110;
        tomato_soup_dim[7][7] = 16'b01100_010100_00110;
        tomato_soup_dim[7][8] = 16'b01100_010101_00111;
        tomato_soup_dim[7][9] = 16'b01100_010101_00111;
        tomato_soup_dim[7][10] = 16'b01100_010101_00111;
        tomato_soup_dim[7][11] = 16'b01100_010101_00111;
        tomato_soup_dim[7][12] = 16'b01100_010101_00110;
        tomato_soup_dim[7][13] = 16'b01100_010101_00111;
        tomato_soup_dim[7][14] = 16'b01100_010101_00111;
        tomato_soup_dim[7][15] = 16'b01100_010101_00110;
        tomato_soup_dim[7][16] = 16'b01100_010101_00111;
        tomato_soup_dim[7][17] = 16'b01101_010101_00111;
        tomato_soup_dim[7][18] = 16'b01100_010100_00110;
        tomato_soup_dim[7][19] = 16'b01100_010101_00110;
        tomato_soup_dim[7][20] = 16'b01101_010110_00111;
        tomato_soup_dim[7][21] = 16'b01101_010101_00111;
        tomato_soup_dim[7][22] = 16'b01100_010101_00111;
        tomato_soup_dim[7][23] = 16'b01101_010101_00111;
        tomato_soup_dim[7][24] = 16'b01100_010101_00110;
        tomato_soup_dim[7][25] = 16'b01011_011111_01010;
        tomato_soup_dim[7][26] = 16'b01011_011111_01010;
        tomato_soup_dim[7][27] = 16'b01011_011111_01010;
        tomato_soup_dim[7][28] = 16'b01011_011111_01010;
        tomato_soup_dim[7][29] = 16'b01011_011111_01010;
        tomato_soup_dim[7][30] = 16'b01011_011111_01010;
        tomato_soup_dim[7][31] = 16'b01011_011111_01010;
        tomato_soup_dim[8][0] = 16'b01011_011111_01010;
        tomato_soup_dim[8][1] = 16'b01011_011111_01010;
        tomato_soup_dim[8][2] = 16'b01011_011111_01010;
        tomato_soup_dim[8][3] = 16'b01011_011111_01010;
        tomato_soup_dim[8][4] = 16'b01011_011111_01010;
        tomato_soup_dim[8][5] = 16'b01100_010100_00110;
        tomato_soup_dim[8][6] = 16'b01100_010100_00110;
        tomato_soup_dim[8][7] = 16'b01100_010101_00111;
        tomato_soup_dim[8][8] = 16'b01100_010101_00111;
        tomato_soup_dim[8][9] = 16'b01100_010100_00110;
        tomato_soup_dim[8][10] = 16'b01100_010101_00111;
        tomato_soup_dim[8][11] = 16'b01100_010101_00110;
        tomato_soup_dim[8][12] = 16'b01100_010100_00110;
        tomato_soup_dim[8][13] = 16'b01100_010100_00110;
        tomato_soup_dim[8][14] = 16'b01100_010100_00110;
        tomato_soup_dim[8][15] = 16'b01100_010101_00111;
        tomato_soup_dim[8][16] = 16'b01100_010100_00110;
        tomato_soup_dim[8][17] = 16'b01100_010100_00110;
        tomato_soup_dim[8][18] = 16'b01100_010100_00110;
        tomato_soup_dim[8][19] = 16'b01100_010100_00110;
        tomato_soup_dim[8][20] = 16'b01100_010101_00111;
        tomato_soup_dim[8][21] = 16'b01100_010100_00110;
        tomato_soup_dim[8][22] = 16'b01100_010101_00111;
        tomato_soup_dim[8][23] = 16'b01100_010101_00111;
        tomato_soup_dim[8][24] = 16'b01100_010101_00111;
        tomato_soup_dim[8][25] = 16'b01100_010101_00110;
        tomato_soup_dim[8][26] = 16'b01011_011111_01010;
        tomato_soup_dim[8][27] = 16'b01011_011111_01010;
        tomato_soup_dim[8][28] = 16'b01011_011111_01010;
        tomato_soup_dim[8][29] = 16'b01011_011111_01010;
        tomato_soup_dim[8][30] = 16'b01011_011111_01010;
        tomato_soup_dim[8][31] = 16'b01011_011111_01010;
        tomato_soup_dim[9][0] = 16'b01011_011111_01010;
        tomato_soup_dim[9][1] = 16'b01011_011111_01010;
        tomato_soup_dim[9][2] = 16'b01011_011111_01010;
        tomato_soup_dim[9][3] = 16'b01011_011111_01010;
        tomato_soup_dim[9][4] = 16'b01011_011111_01010;
        tomato_soup_dim[9][5] = 16'b01100_010101_00110;
        tomato_soup_dim[9][6] = 16'b01100_010101_00111;
        tomato_soup_dim[9][7] = 16'b01100_010100_00110;
        tomato_soup_dim[9][8] = 16'b01100_010100_00110;
        tomato_soup_dim[9][9] = 16'b01100_010101_00111;
        tomato_soup_dim[9][10] = 16'b01100_010101_00111;
        tomato_soup_dim[9][11] = 16'b01100_010101_00111;
        tomato_soup_dim[9][12] = 16'b01101_010110_01000;
        tomato_soup_dim[9][13] = 16'b01101_010111_01000;
        tomato_soup_dim[9][14] = 16'b01101_010110_01000;
        tomato_soup_dim[9][15] = 16'b01101_010110_00111;
        tomato_soup_dim[9][16] = 16'b01101_010110_01000;
        tomato_soup_dim[9][17] = 16'b01101_010111_01000;
        tomato_soup_dim[9][18] = 16'b01101_010111_01000;
        tomato_soup_dim[9][19] = 16'b01101_010110_01000;
        tomato_soup_dim[9][20] = 16'b01100_010101_00110;
        tomato_soup_dim[9][21] = 16'b01100_010100_00110;
        tomato_soup_dim[9][22] = 16'b01100_010101_00110;
        tomato_soup_dim[9][23] = 16'b01100_010101_00110;
        tomato_soup_dim[9][24] = 16'b01100_010101_00111;
        tomato_soup_dim[9][25] = 16'b01100_010100_00110;
        tomato_soup_dim[9][26] = 16'b01100_010100_00110;
        tomato_soup_dim[9][27] = 16'b01011_011111_01010;
        tomato_soup_dim[9][28] = 16'b01011_011111_01010;
        tomato_soup_dim[9][29] = 16'b01011_011111_01010;
        tomato_soup_dim[9][30] = 16'b01011_011111_01010;
        tomato_soup_dim[9][31] = 16'b01011_011111_01010;
        tomato_soup_dim[10][0] = 16'b01011_011111_01010;
        tomato_soup_dim[10][1] = 16'b01011_011111_01010;
        tomato_soup_dim[10][2] = 16'b01011_011111_01010;
        tomato_soup_dim[10][3] = 16'b01011_011111_01010;
        tomato_soup_dim[10][4] = 16'b01100_010100_00110;
        tomato_soup_dim[10][5] = 16'b01100_010100_00110;
        tomato_soup_dim[10][6] = 16'b01100_010100_00110;
        tomato_soup_dim[10][7] = 16'b01100_010100_00110;
        tomato_soup_dim[10][8] = 16'b01101_010110_01000;
        tomato_soup_dim[10][9] = 16'b01101_010111_01000;
        tomato_soup_dim[10][10] = 16'b01101_010111_01000;
        tomato_soup_dim[10][11] = 16'b01101_010110_00111;
        tomato_soup_dim[10][12] = 16'b01100_010100_00110;
        tomato_soup_dim[10][13] = 16'b01100_001111_00011;
        tomato_soup_dim[10][14] = 16'b01100_001100_00010;
        tomato_soup_dim[10][15] = 16'b01100_001100_00010;
        tomato_soup_dim[10][16] = 16'b01100_001101_00011;
        tomato_soup_dim[10][17] = 16'b01100_001110_00011;
        tomato_soup_dim[10][18] = 16'b01100_010001_00101;
        tomato_soup_dim[10][19] = 16'b01101_010110_00111;
        tomato_soup_dim[10][20] = 16'b01101_010110_00111;
        tomato_soup_dim[10][21] = 16'b01101_010110_00111;
        tomato_soup_dim[10][22] = 16'b01101_010110_01000;
        tomato_soup_dim[10][23] = 16'b01100_010101_00110;
        tomato_soup_dim[10][24] = 16'b01100_010100_00110;
        tomato_soup_dim[10][25] = 16'b01100_010101_00110;
        tomato_soup_dim[10][26] = 16'b01100_010101_00110;
        tomato_soup_dim[10][27] = 16'b01011_011111_01010;
        tomato_soup_dim[10][28] = 16'b01011_011111_01010;
        tomato_soup_dim[10][29] = 16'b01011_011111_01010;
        tomato_soup_dim[10][30] = 16'b01011_011111_01010;
        tomato_soup_dim[10][31] = 16'b01011_011111_01010;
        tomato_soup_dim[11][0] = 16'b01011_011111_01010;
        tomato_soup_dim[11][1] = 16'b01011_011111_01010;
        tomato_soup_dim[11][2] = 16'b01011_011111_01010;
        tomato_soup_dim[11][3] = 16'b01011_011111_01010;
        tomato_soup_dim[11][4] = 16'b01100_010100_00110;
        tomato_soup_dim[11][5] = 16'b01100_010100_00110;
        tomato_soup_dim[11][6] = 16'b01101_010110_01000;
        tomato_soup_dim[11][7] = 16'b01101_010110_01000;
        tomato_soup_dim[11][8] = 16'b01101_010110_01000;
        tomato_soup_dim[11][9] = 16'b01100_001110_00011;
        tomato_soup_dim[11][10] = 16'b01011_001001_00001;
        tomato_soup_dim[11][11] = 16'b01011_000110_00000;
        tomato_soup_dim[11][12] = 16'b01011_000110_00000;
        tomato_soup_dim[11][13] = 16'b01011_000101_00000;
        tomato_soup_dim[11][14] = 16'b01100_000110_00000;
        tomato_soup_dim[11][15] = 16'b01011_000110_00000;
        tomato_soup_dim[11][16] = 16'b01011_000110_00000;
        tomato_soup_dim[11][17] = 16'b01011_000101_00000;
        tomato_soup_dim[11][18] = 16'b01011_000110_00000;
        tomato_soup_dim[11][19] = 16'b01011_000101_00000;
        tomato_soup_dim[11][20] = 16'b01011_000101_00000;
        tomato_soup_dim[11][21] = 16'b01100_001100_00010;
        tomato_soup_dim[11][22] = 16'b01101_010111_01000;
        tomato_soup_dim[11][23] = 16'b01101_011000_01001;
        tomato_soup_dim[11][24] = 16'b01101_010111_01000;
        tomato_soup_dim[11][25] = 16'b01100_010100_00110;
        tomato_soup_dim[11][26] = 16'b01100_010100_00110;
        tomato_soup_dim[11][27] = 16'b01100_010100_00110;
        tomato_soup_dim[11][28] = 16'b01011_011111_01010;
        tomato_soup_dim[11][29] = 16'b01011_011111_01010;
        tomato_soup_dim[11][30] = 16'b01011_011111_01010;
        tomato_soup_dim[11][31] = 16'b01011_011111_01010;
        tomato_soup_dim[12][0] = 16'b01011_011111_01010;
        tomato_soup_dim[12][1] = 16'b01011_011111_01010;
        tomato_soup_dim[12][2] = 16'b01011_011111_01010;
        tomato_soup_dim[12][3] = 16'b01100_010100_00110;
        tomato_soup_dim[12][4] = 16'b01100_010100_00110;
        tomato_soup_dim[12][5] = 16'b01101_010111_01000;
        tomato_soup_dim[12][6] = 16'b01101_010101_00111;
        tomato_soup_dim[12][7] = 16'b01100_001011_00010;
        tomato_soup_dim[12][8] = 16'b01011_000101_00000;
        tomato_soup_dim[12][9] = 16'b01011_000101_00000;
        tomato_soup_dim[12][10] = 16'b01011_000101_00000;
        tomato_soup_dim[12][11] = 16'b01011_000110_00000;
        tomato_soup_dim[12][12] = 16'b01011_000110_00000;
        tomato_soup_dim[12][13] = 16'b01011_000110_00000;
        tomato_soup_dim[12][14] = 16'b01100_000111_00000;
        tomato_soup_dim[12][15] = 16'b01100_000111_00000;
        tomato_soup_dim[12][16] = 16'b01100_000111_00000;
        tomato_soup_dim[12][17] = 16'b01100_000110_00000;
        tomato_soup_dim[12][18] = 16'b01100_000111_00000;
        tomato_soup_dim[12][19] = 16'b01100_000110_00000;
        tomato_soup_dim[12][20] = 16'b01100_000110_00000;
        tomato_soup_dim[12][21] = 16'b01100_000111_00000;
        tomato_soup_dim[12][22] = 16'b01011_000110_00000;
        tomato_soup_dim[12][23] = 16'b01100_001011_00010;
        tomato_soup_dim[12][24] = 16'b01101_010101_00111;
        tomato_soup_dim[12][25] = 16'b01101_011000_01001;
        tomato_soup_dim[12][26] = 16'b01100_010100_00110;
        tomato_soup_dim[12][27] = 16'b01100_010100_00110;
        tomato_soup_dim[12][28] = 16'b01011_011111_01010;
        tomato_soup_dim[12][29] = 16'b01011_011111_01010;
        tomato_soup_dim[12][30] = 16'b01011_011111_01010;
        tomato_soup_dim[12][31] = 16'b01011_011111_01010;
        tomato_soup_dim[13][0] = 16'b01011_011111_01010;
        tomato_soup_dim[13][1] = 16'b01011_011111_01010;
        tomato_soup_dim[13][2] = 16'b01011_011111_01010;
        tomato_soup_dim[13][3] = 16'b01100_010100_00110;
        tomato_soup_dim[13][4] = 16'b01101_010110_00111;
        tomato_soup_dim[13][5] = 16'b01100_001111_00100;
        tomato_soup_dim[13][6] = 16'b01011_000110_00000;
        tomato_soup_dim[13][7] = 16'b01011_000101_00000;
        tomato_soup_dim[13][8] = 16'b01011_000110_00000;
        tomato_soup_dim[13][9] = 16'b01011_000101_00000;
        tomato_soup_dim[13][10] = 16'b01100_000111_00000;
        tomato_soup_dim[13][11] = 16'b01100_000111_00000;
        tomato_soup_dim[13][12] = 16'b01100_000111_00000;
        tomato_soup_dim[13][13] = 16'b01100_000111_00000;
        tomato_soup_dim[13][14] = 16'b01100_000111_00000;
        tomato_soup_dim[13][15] = 16'b01100_000111_00000;
        tomato_soup_dim[13][16] = 16'b01100_000111_00000;
        tomato_soup_dim[13][17] = 16'b01100_000111_00000;
        tomato_soup_dim[13][18] = 16'b01100_000111_00001;
        tomato_soup_dim[13][19] = 16'b01100_000111_00000;
        tomato_soup_dim[13][20] = 16'b01100_000111_00000;
        tomato_soup_dim[13][21] = 16'b01100_000111_00000;
        tomato_soup_dim[13][22] = 16'b01100_000111_00000;
        tomato_soup_dim[13][23] = 16'b01100_000111_00000;
        tomato_soup_dim[13][24] = 16'b01100_000110_00000;
        tomato_soup_dim[13][25] = 16'b01100_010001_00101;
        tomato_soup_dim[13][26] = 16'b01110_011000_01001;
        tomato_soup_dim[13][27] = 16'b01100_010101_00110;
        tomato_soup_dim[13][28] = 16'b01100_010100_00110;
        tomato_soup_dim[13][29] = 16'b01011_011111_01010;
        tomato_soup_dim[13][30] = 16'b01011_011111_01010;
        tomato_soup_dim[13][31] = 16'b01011_011111_01010;
        tomato_soup_dim[14][0] = 16'b01011_011111_01010;
        tomato_soup_dim[14][1] = 16'b01011_011111_01010;
        tomato_soup_dim[14][2] = 16'b01101_010111_01000;
        tomato_soup_dim[14][3] = 16'b01101_010111_01000;
        tomato_soup_dim[14][4] = 16'b01100_010001_00100;
        tomato_soup_dim[14][5] = 16'b01011_000101_00000;
        tomato_soup_dim[14][6] = 16'b01011_000110_00000;
        tomato_soup_dim[14][7] = 16'b01011_000110_00000;
        tomato_soup_dim[14][8] = 16'b01100_000111_00000;
        tomato_soup_dim[14][9] = 16'b01100_000111_00001;
        tomato_soup_dim[14][10] = 16'b01100_000110_00000;
        tomato_soup_dim[14][11] = 16'b01100_000111_00001;
        tomato_soup_dim[14][12] = 16'b01100_000111_00000;
        tomato_soup_dim[14][13] = 16'b01100_000110_00000;
        tomato_soup_dim[14][14] = 16'b01100_000111_00000;
        tomato_soup_dim[14][15] = 16'b01100_000110_00000;
        tomato_soup_dim[14][16] = 16'b01011_000110_00000;
        tomato_soup_dim[14][17] = 16'b01100_000110_00000;
        tomato_soup_dim[14][18] = 16'b01011_000110_00000;
        tomato_soup_dim[14][19] = 16'b01011_000110_00000;
        tomato_soup_dim[14][20] = 16'b01011_000110_00000;
        tomato_soup_dim[14][21] = 16'b01011_000110_00000;
        tomato_soup_dim[14][22] = 16'b01100_000111_00000;
        tomato_soup_dim[14][23] = 16'b01100_000111_00001;
        tomato_soup_dim[14][24] = 16'b01100_000111_00000;
        tomato_soup_dim[14][25] = 16'b01100_000111_00000;
        tomato_soup_dim[14][26] = 16'b01100_001101_00011;
        tomato_soup_dim[14][27] = 16'b01101_011000_01001;
        tomato_soup_dim[14][28] = 16'b01100_010100_00110;
        tomato_soup_dim[14][29] = 16'b01011_011111_01010;
        tomato_soup_dim[14][30] = 16'b01011_011111_01010;
        tomato_soup_dim[14][31] = 16'b01011_011111_01010;
        tomato_soup_dim[15][0] = 16'b01011_011111_01010;
        tomato_soup_dim[15][1] = 16'b01011_011111_01010;
        tomato_soup_dim[15][2] = 16'b01110_011001_01001;
        tomato_soup_dim[15][3] = 16'b01110_011000_01001;
        tomato_soup_dim[15][4] = 16'b01011_000110_00000;
        tomato_soup_dim[15][5] = 16'b01011_000101_00000;
        tomato_soup_dim[15][6] = 16'b01011_000110_00000;
        tomato_soup_dim[15][7] = 16'b01100_000110_00000;
        tomato_soup_dim[15][8] = 16'b01100_000111_00000;
        tomato_soup_dim[15][9] = 16'b01101_001000_00001;
        tomato_soup_dim[15][10] = 16'b01100_000111_00000;
        tomato_soup_dim[15][11] = 16'b01100_000110_00000;
        tomato_soup_dim[15][12] = 16'b01100_000111_00000;
        tomato_soup_dim[15][13] = 16'b01011_000110_00000;
        tomato_soup_dim[15][14] = 16'b01100_000110_00000;
        tomato_soup_dim[15][15] = 16'b01100_000110_00000;
        tomato_soup_dim[15][16] = 16'b01100_000111_00000;
        tomato_soup_dim[15][17] = 16'b01100_000111_00000;
        tomato_soup_dim[15][18] = 16'b01100_000111_00000;
        tomato_soup_dim[15][19] = 16'b01100_000110_00000;
        tomato_soup_dim[15][20] = 16'b01011_000110_00000;
        tomato_soup_dim[15][21] = 16'b01011_000110_00000;
        tomato_soup_dim[15][22] = 16'b01011_000110_00000;
        tomato_soup_dim[15][23] = 16'b01100_000111_00000;
        tomato_soup_dim[15][24] = 16'b01100_000111_00000;
        tomato_soup_dim[15][25] = 16'b01100_000111_00000;
        tomato_soup_dim[15][26] = 16'b01011_000101_00000;
        tomato_soup_dim[15][27] = 16'b01100_010010_00101;
        tomato_soup_dim[15][28] = 16'b01101_010111_01000;
        tomato_soup_dim[15][29] = 16'b01011_011111_01010;
        tomato_soup_dim[15][30] = 16'b01011_011111_01010;
        tomato_soup_dim[15][31] = 16'b01011_011111_01010;
        tomato_soup_dim[16][0] = 16'b01011_011111_01010;
        tomato_soup_dim[16][1] = 16'b01011_011111_01010;
        tomato_soup_dim[16][2] = 16'b01101_011000_01001;
        tomato_soup_dim[16][3] = 16'b01101_011000_01001;
        tomato_soup_dim[16][4] = 16'b01011_000101_00000;
        tomato_soup_dim[16][5] = 16'b01011_000101_00000;
        tomato_soup_dim[16][6] = 16'b01011_000110_00000;
        tomato_soup_dim[16][7] = 16'b01100_000111_00001;
        tomato_soup_dim[16][8] = 16'b01100_000111_00001;
        tomato_soup_dim[16][9] = 16'b01100_000111_00001;
        tomato_soup_dim[16][10] = 16'b01100_000110_00000;
        tomato_soup_dim[16][11] = 16'b01100_000111_00000;
        tomato_soup_dim[16][12] = 16'b01100_000111_00001;
        tomato_soup_dim[16][13] = 16'b01100_000110_00000;
        tomato_soup_dim[16][14] = 16'b01100_000111_00001;
        tomato_soup_dim[16][15] = 16'b01100_000111_00000;
        tomato_soup_dim[16][16] = 16'b01100_000111_00000;
        tomato_soup_dim[16][17] = 16'b01100_000111_00001;
        tomato_soup_dim[16][18] = 16'b01100_000111_00001;
        tomato_soup_dim[16][19] = 16'b01100_000110_00000;
        tomato_soup_dim[16][20] = 16'b01011_000110_00000;
        tomato_soup_dim[16][21] = 16'b00110_001101_00001;
        tomato_soup_dim[16][22] = 16'b00110_001101_00001;
        tomato_soup_dim[16][23] = 16'b01011_000110_00000;
        tomato_soup_dim[16][24] = 16'b01100_000110_00000;
        tomato_soup_dim[16][25] = 16'b01100_000111_00001;
        tomato_soup_dim[16][26] = 16'b01011_000101_00000;
        tomato_soup_dim[16][27] = 16'b01011_001001_00001;
        tomato_soup_dim[16][28] = 16'b01101_011000_01001;
        tomato_soup_dim[16][29] = 16'b01011_011111_01010;
        tomato_soup_dim[16][30] = 16'b01011_011111_01010;
        tomato_soup_dim[16][31] = 16'b01011_011111_01010;
        tomato_soup_dim[17][0] = 16'b01011_011111_01010;
        tomato_soup_dim[17][1] = 16'b01011_011111_01010;
        tomato_soup_dim[17][2] = 16'b01110_011001_01010;
        tomato_soup_dim[17][3] = 16'b01101_010110_00111;
        tomato_soup_dim[17][4] = 16'b01011_000111_00001;
        tomato_soup_dim[17][5] = 16'b01011_000101_00000;
        tomato_soup_dim[17][6] = 16'b01011_000110_00000;
        tomato_soup_dim[17][7] = 16'b01011_000110_00000;
        tomato_soup_dim[17][8] = 16'b01100_000111_00001;
        tomato_soup_dim[17][9] = 16'b01100_000111_00001;
        tomato_soup_dim[17][10] = 16'b01100_000110_00000;
        tomato_soup_dim[17][11] = 16'b01100_000110_00000;
        tomato_soup_dim[17][12] = 16'b01100_000111_00001;
        tomato_soup_dim[17][13] = 16'b01100_000110_00000;
        tomato_soup_dim[17][14] = 16'b01100_000111_00000;
        tomato_soup_dim[17][15] = 16'b01100_000111_00001;
        tomato_soup_dim[17][16] = 16'b01100_000111_00001;
        tomato_soup_dim[17][17] = 16'b01100_000111_00000;
        tomato_soup_dim[17][18] = 16'b01100_000111_00000;
        tomato_soup_dim[17][19] = 16'b00110_001101_00001;
        tomato_soup_dim[17][20] = 16'b00110_001100_00001;
        tomato_soup_dim[17][21] = 16'b00110_001101_00001;
        tomato_soup_dim[17][22] = 16'b00101_001100_00001;
        tomato_soup_dim[17][23] = 16'b00101_001011_00001;
        tomato_soup_dim[17][24] = 16'b01011_000110_00000;
        tomato_soup_dim[17][25] = 16'b01100_001000_00001;
        tomato_soup_dim[17][26] = 16'b01011_000101_00000;
        tomato_soup_dim[17][27] = 16'b01011_001010_00010;
        tomato_soup_dim[17][28] = 16'b01110_011001_01001;
        tomato_soup_dim[17][29] = 16'b01011_011111_01010;
        tomato_soup_dim[17][30] = 16'b01011_011111_01010;
        tomato_soup_dim[17][31] = 16'b01011_011111_01010;
        tomato_soup_dim[18][0] = 16'b01011_011111_01010;
        tomato_soup_dim[18][1] = 16'b01011_011111_01010;
        tomato_soup_dim[18][2] = 16'b01110_011001_01010;
        tomato_soup_dim[18][3] = 16'b01101_010101_00111;
        tomato_soup_dim[18][4] = 16'b01100_001110_00011;
        tomato_soup_dim[18][5] = 16'b01011_000110_00000;
        tomato_soup_dim[18][6] = 16'b01011_000101_00000;
        tomato_soup_dim[18][7] = 16'b01011_000110_00000;
        tomato_soup_dim[18][8] = 16'b01100_000111_00001;
        tomato_soup_dim[18][9] = 16'b01100_000111_00000;
        tomato_soup_dim[18][10] = 16'b01100_000111_00001;
        tomato_soup_dim[18][11] = 16'b01100_000110_00000;
        tomato_soup_dim[18][12] = 16'b01100_000110_00000;
        tomato_soup_dim[18][13] = 16'b01011_000110_00000;
        tomato_soup_dim[18][14] = 16'b01100_000110_00000;
        tomato_soup_dim[18][15] = 16'b01100_000110_00000;
        tomato_soup_dim[18][16] = 16'b01100_000111_00000;
        tomato_soup_dim[18][17] = 16'b01100_000110_00000;
        tomato_soup_dim[18][18] = 16'b00110_001101_00001;
        tomato_soup_dim[18][19] = 16'b00110_001101_00001;
        tomato_soup_dim[18][20] = 16'b00101_001100_00001;
        tomato_soup_dim[18][21] = 16'b00110_001110_00001;
        tomato_soup_dim[18][22] = 16'b00110_001110_00001;
        tomato_soup_dim[18][23] = 16'b00110_001101_00001;
        tomato_soup_dim[18][24] = 16'b01011_000110_00000;
        tomato_soup_dim[18][25] = 16'b01100_000110_00000;
        tomato_soup_dim[18][26] = 16'b01011_000101_00000;
        tomato_soup_dim[18][27] = 16'b01100_010100_00110;
        tomato_soup_dim[18][28] = 16'b01110_011001_01010;
        tomato_soup_dim[18][29] = 16'b01011_011111_01010;
        tomato_soup_dim[18][30] = 16'b01011_011111_01010;
        tomato_soup_dim[18][31] = 16'b01011_011111_01010;
        tomato_soup_dim[19][0] = 16'b01011_011111_01010;
        tomato_soup_dim[19][1] = 16'b01011_011111_01010;
        tomato_soup_dim[19][2] = 16'b01011_011111_01010;
        tomato_soup_dim[19][3] = 16'b01101_010111_01000;
        tomato_soup_dim[19][4] = 16'b01100_010100_00110;
        tomato_soup_dim[19][5] = 16'b01011_001100_00010;
        tomato_soup_dim[19][6] = 16'b01011_000110_00000;
        tomato_soup_dim[19][7] = 16'b01011_000101_00000;
        tomato_soup_dim[19][8] = 16'b01100_000111_00001;
        tomato_soup_dim[19][9] = 16'b01100_000111_00000;
        tomato_soup_dim[19][10] = 16'b01100_000111_00001;
        tomato_soup_dim[19][11] = 16'b01100_000111_00000;
        tomato_soup_dim[19][12] = 16'b01100_000111_00000;
        tomato_soup_dim[19][13] = 16'b01100_000110_00000;
        tomato_soup_dim[19][14] = 16'b01100_000110_00000;
        tomato_soup_dim[19][15] = 16'b01100_000110_00000;
        tomato_soup_dim[19][16] = 16'b01100_000110_00000;
        tomato_soup_dim[19][17] = 16'b01100_000110_00000;
        tomato_soup_dim[19][18] = 16'b00110_001101_00001;
        tomato_soup_dim[19][19] = 16'b00110_001100_00001;
        tomato_soup_dim[19][20] = 16'b00101_001100_00001;
        tomato_soup_dim[19][21] = 16'b00101_001011_00001;
        tomato_soup_dim[19][22] = 16'b00101_001010_00001;
        tomato_soup_dim[19][23] = 16'b01011_000101_00000;
        tomato_soup_dim[19][24] = 16'b01011_000110_00000;
        tomato_soup_dim[19][25] = 16'b01011_000110_00000;
        tomato_soup_dim[19][26] = 16'b01100_010000_00100;
        tomato_soup_dim[19][27] = 16'b01101_010110_00111;
        tomato_soup_dim[19][28] = 16'b01110_011001_01010;
        tomato_soup_dim[19][29] = 16'b01011_011111_01010;
        tomato_soup_dim[19][30] = 16'b01011_011111_01010;
        tomato_soup_dim[19][31] = 16'b01011_011111_01010;
        tomato_soup_dim[20][0] = 16'b01011_011111_01010;
        tomato_soup_dim[20][1] = 16'b01011_011111_01010;
        tomato_soup_dim[20][2] = 16'b01011_011111_01010;
        tomato_soup_dim[20][3] = 16'b01101_010110_00111;
        tomato_soup_dim[20][4] = 16'b01101_010101_00111;
        tomato_soup_dim[20][5] = 16'b01100_010101_00111;
        tomato_soup_dim[20][6] = 16'b01100_001111_00011;
        tomato_soup_dim[20][7] = 16'b01011_000110_00000;
        tomato_soup_dim[20][8] = 16'b01011_000101_00000;
        tomato_soup_dim[20][9] = 16'b01011_000101_00000;
        tomato_soup_dim[20][10] = 16'b01100_000111_00001;
        tomato_soup_dim[20][11] = 16'b01100_000111_00001;
        tomato_soup_dim[20][12] = 16'b01100_000111_00000;
        tomato_soup_dim[20][13] = 16'b01100_000110_00000;
        tomato_soup_dim[20][14] = 16'b01100_000111_00000;
        tomato_soup_dim[20][15] = 16'b01100_000111_00000;
        tomato_soup_dim[20][16] = 16'b01100_000111_00001;
        tomato_soup_dim[20][17] = 16'b01100_000111_00000;
        tomato_soup_dim[20][18] = 16'b01100_000111_00000;
        tomato_soup_dim[20][19] = 16'b00110_001101_00001;
        tomato_soup_dim[20][20] = 16'b00110_001101_00001;
        tomato_soup_dim[20][21] = 16'b01011_000101_00000;
        tomato_soup_dim[20][22] = 16'b01011_000101_00000;
        tomato_soup_dim[20][23] = 16'b01011_000110_00000;
        tomato_soup_dim[20][24] = 16'b01011_000110_00000;
        tomato_soup_dim[20][25] = 16'b01100_010000_00100;
        tomato_soup_dim[20][26] = 16'b01101_010101_00111;
        tomato_soup_dim[20][27] = 16'b01101_010111_01000;
        tomato_soup_dim[20][28] = 16'b01101_011000_01001;
        tomato_soup_dim[20][29] = 16'b01011_011111_01010;
        tomato_soup_dim[20][30] = 16'b01011_011111_01010;
        tomato_soup_dim[20][31] = 16'b01011_011111_01010;
        tomato_soup_dim[21][0] = 16'b01011_011111_01010;
        tomato_soup_dim[21][1] = 16'b01011_011111_01010;
        tomato_soup_dim[21][2] = 16'b01011_011111_01010;
        tomato_soup_dim[21][3] = 16'b01011_011111_01010;
        tomato_soup_dim[21][4] = 16'b01101_010111_01000;
        tomato_soup_dim[21][5] = 16'b01100_010101_00111;
        tomato_soup_dim[21][6] = 16'b01100_010100_00110;
        tomato_soup_dim[21][7] = 16'b01100_010100_00110;
        tomato_soup_dim[21][8] = 16'b01011_001010_00001;
        tomato_soup_dim[21][9] = 16'b01011_000110_00000;
        tomato_soup_dim[21][10] = 16'b01011_000110_00000;
        tomato_soup_dim[21][11] = 16'b01011_000101_00000;
        tomato_soup_dim[21][12] = 16'b01011_000101_00000;
        tomato_soup_dim[21][13] = 16'b01011_000101_00000;
        tomato_soup_dim[21][14] = 16'b01011_000110_00000;
        tomato_soup_dim[21][15] = 16'b01100_000111_00000;
        tomato_soup_dim[21][16] = 16'b01100_000111_00000;
        tomato_soup_dim[21][17] = 16'b01100_000111_00000;
        tomato_soup_dim[21][18] = 16'b01100_000111_00000;
        tomato_soup_dim[21][19] = 16'b01100_000110_00000;
        tomato_soup_dim[21][20] = 16'b01011_000110_00000;
        tomato_soup_dim[21][21] = 16'b01011_000110_00000;
        tomato_soup_dim[21][22] = 16'b01011_000110_00000;
        tomato_soup_dim[21][23] = 16'b01100_001011_00010;
        tomato_soup_dim[21][24] = 16'b01100_010100_00110;
        tomato_soup_dim[21][25] = 16'b01100_010100_00110;
        tomato_soup_dim[21][26] = 16'b01101_010101_00111;
        tomato_soup_dim[21][27] = 16'b01101_011000_01001;
        tomato_soup_dim[21][28] = 16'b01011_011111_01010;
        tomato_soup_dim[21][29] = 16'b01011_011111_01010;
        tomato_soup_dim[21][30] = 16'b01011_011111_01010;
        tomato_soup_dim[21][31] = 16'b01011_011111_01010;
        tomato_soup_dim[22][0] = 16'b01011_011111_01010;
        tomato_soup_dim[22][1] = 16'b01011_011111_01010;
        tomato_soup_dim[22][2] = 16'b01011_011111_01010;
        tomato_soup_dim[22][3] = 16'b01011_011111_01010;
        tomato_soup_dim[22][4] = 16'b01011_011111_01010;
        tomato_soup_dim[22][5] = 16'b01101_011000_01001;
        tomato_soup_dim[22][6] = 16'b01100_010101_00110;
        tomato_soup_dim[22][7] = 16'b01100_010100_00110;
        tomato_soup_dim[22][8] = 16'b01100_010100_00110;
        tomato_soup_dim[22][9] = 16'b01100_010100_00110;
        tomato_soup_dim[22][10] = 16'b01100_010100_00110;
        tomato_soup_dim[22][11] = 16'b01100_001010_00001;
        tomato_soup_dim[22][12] = 16'b01011_000110_00000;
        tomato_soup_dim[22][13] = 16'b01011_000101_00000;
        tomato_soup_dim[22][14] = 16'b01011_000110_00000;
        tomato_soup_dim[22][15] = 16'b01011_000110_00000;
        tomato_soup_dim[22][16] = 16'b01011_000110_00000;
        tomato_soup_dim[22][17] = 16'b01100_000111_00000;
        tomato_soup_dim[22][18] = 16'b01100_000111_00000;
        tomato_soup_dim[22][19] = 16'b01100_000110_00000;
        tomato_soup_dim[22][20] = 16'b01100_001011_00010;
        tomato_soup_dim[22][21] = 16'b01100_010100_00110;
        tomato_soup_dim[22][22] = 16'b01100_010100_00110;
        tomato_soup_dim[22][23] = 16'b01100_010100_00110;
        tomato_soup_dim[22][24] = 16'b01100_010100_00110;
        tomato_soup_dim[22][25] = 16'b01100_010101_00111;
        tomato_soup_dim[22][26] = 16'b01101_010111_01000;
        tomato_soup_dim[22][27] = 16'b01011_011111_01010;
        tomato_soup_dim[22][28] = 16'b01011_011111_01010;
        tomato_soup_dim[22][29] = 16'b01011_011111_01010;
        tomato_soup_dim[22][30] = 16'b01011_011111_01010;
        tomato_soup_dim[22][31] = 16'b01011_011111_01010;
        tomato_soup_dim[23][0] = 16'b01011_011111_01010;
        tomato_soup_dim[23][1] = 16'b01011_011111_01010;
        tomato_soup_dim[23][2] = 16'b01011_011111_01010;
        tomato_soup_dim[23][3] = 16'b01011_011111_01010;
        tomato_soup_dim[23][4] = 16'b01011_011111_01010;
        tomato_soup_dim[23][5] = 16'b01011_011111_01010;
        tomato_soup_dim[23][6] = 16'b01101_010111_01000;
        tomato_soup_dim[23][7] = 16'b01101_010111_01000;
        tomato_soup_dim[23][8] = 16'b01100_010100_00110;
        tomato_soup_dim[23][9] = 16'b01100_010100_00110;
        tomato_soup_dim[23][10] = 16'b01100_010101_00110;
        tomato_soup_dim[23][11] = 16'b01100_010100_00110;
        tomato_soup_dim[23][12] = 16'b01100_010100_00110;
        tomato_soup_dim[23][13] = 16'b01100_010100_00110;
        tomato_soup_dim[23][14] = 16'b01100_010100_00110;
        tomato_soup_dim[23][15] = 16'b01100_010100_00110;
        tomato_soup_dim[23][16] = 16'b01100_010100_00110;
        tomato_soup_dim[23][17] = 16'b01100_010100_00110;
        tomato_soup_dim[23][18] = 16'b01100_010100_00110;
        tomato_soup_dim[23][19] = 16'b01100_010100_00110;
        tomato_soup_dim[23][20] = 16'b01100_010100_00110;
        tomato_soup_dim[23][21] = 16'b01100_010100_00110;
        tomato_soup_dim[23][22] = 16'b01100_010100_00110;
        tomato_soup_dim[23][23] = 16'b01101_010110_00111;
        tomato_soup_dim[23][24] = 16'b01101_010111_01000;
        tomato_soup_dim[23][25] = 16'b01101_010111_01000;
        tomato_soup_dim[23][26] = 16'b01011_011111_01010;
        tomato_soup_dim[23][27] = 16'b01011_011111_01010;
        tomato_soup_dim[23][28] = 16'b01011_011111_01010;
        tomato_soup_dim[23][29] = 16'b01011_011111_01010;
        tomato_soup_dim[23][30] = 16'b01011_011111_01010;
        tomato_soup_dim[23][31] = 16'b01011_011111_01010;
        tomato_soup_dim[24][0] = 16'b01011_011111_01010;
        tomato_soup_dim[24][1] = 16'b01011_011111_01010;
        tomato_soup_dim[24][2] = 16'b01011_011111_01010;
        tomato_soup_dim[24][3] = 16'b01011_011111_01010;
        tomato_soup_dim[24][4] = 16'b01011_011111_01010;
        tomato_soup_dim[24][5] = 16'b01011_011111_01010;
        tomato_soup_dim[24][6] = 16'b01011_011111_01010;
        tomato_soup_dim[24][7] = 16'b01101_011000_01001;
        tomato_soup_dim[24][8] = 16'b01101_011000_01001;
        tomato_soup_dim[24][9] = 16'b01101_011000_01001;
        tomato_soup_dim[24][10] = 16'b01101_011000_01001;
        tomato_soup_dim[24][11] = 16'b01100_010100_00110;
        tomato_soup_dim[24][12] = 16'b01100_010100_00110;
        tomato_soup_dim[24][13] = 16'b01100_010100_00110;
        tomato_soup_dim[24][14] = 16'b01100_010100_00110;
        tomato_soup_dim[24][15] = 16'b01100_010100_00110;
        tomato_soup_dim[24][16] = 16'b01100_010100_00110;
        tomato_soup_dim[24][17] = 16'b01100_010100_00110;
        tomato_soup_dim[24][18] = 16'b01100_010100_00110;
        tomato_soup_dim[24][19] = 16'b01100_010100_00110;
        tomato_soup_dim[24][20] = 16'b01100_010100_00110;
        tomato_soup_dim[24][21] = 16'b01101_010111_01000;
        tomato_soup_dim[24][22] = 16'b01101_011000_01001;
        tomato_soup_dim[24][23] = 16'b01101_011000_01001;
        tomato_soup_dim[24][24] = 16'b01101_011000_01001;
        tomato_soup_dim[24][25] = 16'b01011_011111_01010;
        tomato_soup_dim[24][26] = 16'b01011_011111_01010;
        tomato_soup_dim[24][27] = 16'b01011_011111_01010;
        tomato_soup_dim[24][28] = 16'b01011_011111_01010;
        tomato_soup_dim[24][29] = 16'b01011_011111_01010;
        tomato_soup_dim[24][30] = 16'b01011_011111_01010;
        tomato_soup_dim[24][31] = 16'b01011_011111_01010;
        tomato_soup_dim[25][0] = 16'b01011_011111_01010;
        tomato_soup_dim[25][1] = 16'b01011_011111_01010;
        tomato_soup_dim[25][2] = 16'b01011_011111_01010;
        tomato_soup_dim[25][3] = 16'b01011_011111_01010;
        tomato_soup_dim[25][4] = 16'b01011_011111_01010;
        tomato_soup_dim[25][5] = 16'b01011_011111_01010;
        tomato_soup_dim[25][6] = 16'b01011_011111_01010;
        tomato_soup_dim[25][7] = 16'b01011_011111_01010;
        tomato_soup_dim[25][8] = 16'b01011_011111_01010;
        tomato_soup_dim[25][9] = 16'b01011_011111_01010;
        tomato_soup_dim[25][10] = 16'b01110_011001_01001;
        tomato_soup_dim[25][11] = 16'b01110_011001_01001;
        tomato_soup_dim[25][12] = 16'b01101_011000_01001;
        tomato_soup_dim[25][13] = 16'b01110_011001_01001;
        tomato_soup_dim[25][14] = 16'b01101_011000_01001;
        tomato_soup_dim[25][15] = 16'b01101_011000_01001;
        tomato_soup_dim[25][16] = 16'b01101_011000_01001;
        tomato_soup_dim[25][17] = 16'b01101_011000_01001;
        tomato_soup_dim[25][18] = 16'b01101_011000_01001;
        tomato_soup_dim[25][19] = 16'b01101_010111_01000;
        tomato_soup_dim[25][20] = 16'b01101_011000_01001;
        tomato_soup_dim[25][21] = 16'b01101_011000_01001;
        tomato_soup_dim[25][22] = 16'b01011_011111_01010;
        tomato_soup_dim[25][23] = 16'b01011_011111_01010;
        tomato_soup_dim[25][24] = 16'b01011_011111_01010;
        tomato_soup_dim[25][25] = 16'b01011_011111_01010;
        tomato_soup_dim[25][26] = 16'b01011_011111_01010;
        tomato_soup_dim[25][27] = 16'b01011_011111_01010;
        tomato_soup_dim[25][28] = 16'b01011_011111_01010;
        tomato_soup_dim[25][29] = 16'b01011_011111_01010;
        tomato_soup_dim[25][30] = 16'b01011_011111_01010;
        tomato_soup_dim[25][31] = 16'b01011_011111_01010;
        tomato_soup_dim[26][0] = 16'b01011_011111_01010;
        tomato_soup_dim[26][1] = 16'b01011_011111_01010;
        tomato_soup_dim[26][2] = 16'b01011_011111_01010;
        tomato_soup_dim[26][3] = 16'b01011_011111_01010;
        tomato_soup_dim[26][4] = 16'b01011_011111_01010;
        tomato_soup_dim[26][5] = 16'b01011_011111_01010;
        tomato_soup_dim[26][6] = 16'b01011_011111_01010;
        tomato_soup_dim[26][7] = 16'b01011_011111_01010;
        tomato_soup_dim[26][8] = 16'b01011_011111_01010;
        tomato_soup_dim[26][9] = 16'b01011_011111_01010;
        tomato_soup_dim[26][10] = 16'b01011_011111_01010;
        tomato_soup_dim[26][11] = 16'b01011_011111_01010;
        tomato_soup_dim[26][12] = 16'b01011_011111_01010;
        tomato_soup_dim[26][13] = 16'b01011_011111_01010;
        tomato_soup_dim[26][14] = 16'b01011_011111_01010;
        tomato_soup_dim[26][15] = 16'b01011_011111_01010;
        tomato_soup_dim[26][16] = 16'b01011_011111_01010;
        tomato_soup_dim[26][17] = 16'b01011_011111_01010;
        tomato_soup_dim[26][18] = 16'b01011_011111_01010;
        tomato_soup_dim[26][19] = 16'b01011_011111_01010;
        tomato_soup_dim[26][20] = 16'b01011_011111_01010;
        tomato_soup_dim[26][21] = 16'b01011_011111_01010;
        tomato_soup_dim[26][22] = 16'b01011_011111_01010;
        tomato_soup_dim[26][23] = 16'b01011_011111_01010;
        tomato_soup_dim[26][24] = 16'b01011_011111_01010;
        tomato_soup_dim[26][25] = 16'b01011_011111_01010;
        tomato_soup_dim[26][26] = 16'b01011_011111_01010;
        tomato_soup_dim[26][27] = 16'b01011_011111_01010;
        tomato_soup_dim[26][28] = 16'b01011_011111_01010;
        tomato_soup_dim[26][29] = 16'b01011_011111_01010;
        tomato_soup_dim[26][30] = 16'b01011_011111_01010;
        tomato_soup_dim[26][31] = 16'b01011_011111_01010;
        tomato_soup_dim[27][0] = 16'b01011_011111_01010;
        tomato_soup_dim[27][1] = 16'b01011_011111_01010;
        tomato_soup_dim[27][2] = 16'b01011_011111_01010;
        tomato_soup_dim[27][3] = 16'b01011_011111_01010;
        tomato_soup_dim[27][4] = 16'b01011_011111_01010;
        tomato_soup_dim[27][5] = 16'b01011_011111_01010;
        tomato_soup_dim[27][6] = 16'b01011_011111_01010;
        tomato_soup_dim[27][7] = 16'b01011_011111_01010;
        tomato_soup_dim[27][8] = 16'b01011_011111_01010;
        tomato_soup_dim[27][9] = 16'b01011_011111_01010;
        tomato_soup_dim[27][10] = 16'b01011_011111_01010;
        tomato_soup_dim[27][11] = 16'b01011_011111_01010;
        tomato_soup_dim[27][12] = 16'b01011_011111_01010;
        tomato_soup_dim[27][13] = 16'b01011_011111_01010;
        tomato_soup_dim[27][14] = 16'b01011_011111_01010;
        tomato_soup_dim[27][15] = 16'b01011_011111_01010;
        tomato_soup_dim[27][16] = 16'b01011_011111_01010;
        tomato_soup_dim[27][17] = 16'b01011_011111_01010;
        tomato_soup_dim[27][18] = 16'b01011_011111_01010;
        tomato_soup_dim[27][19] = 16'b01011_011111_01010;
        tomato_soup_dim[27][20] = 16'b01011_011111_01010;
        tomato_soup_dim[27][21] = 16'b01011_011111_01010;
        tomato_soup_dim[27][22] = 16'b01011_011111_01010;
        tomato_soup_dim[27][23] = 16'b01011_011111_01010;
        tomato_soup_dim[27][24] = 16'b01011_011111_01010;
        tomato_soup_dim[27][25] = 16'b01011_011111_01010;
        tomato_soup_dim[27][26] = 16'b01011_011111_01010;
        tomato_soup_dim[27][27] = 16'b01011_011111_01010;
        tomato_soup_dim[27][28] = 16'b01011_011111_01010;
        tomato_soup_dim[27][29] = 16'b01011_011111_01010;
        tomato_soup_dim[27][30] = 16'b01011_011111_01010;
        tomato_soup_dim[27][31] = 16'b01011_011111_01010;
        tomato_soup_dim[28][0] = 16'b01011_011111_01010;
        tomato_soup_dim[28][1] = 16'b01011_011111_01010;
        tomato_soup_dim[28][2] = 16'b01011_011111_01010;
        tomato_soup_dim[28][3] = 16'b01011_011111_01010;
        tomato_soup_dim[28][4] = 16'b01011_011111_01010;
        tomato_soup_dim[28][5] = 16'b01011_011111_01010;
        tomato_soup_dim[28][6] = 16'b01011_011111_01010;
        tomato_soup_dim[28][7] = 16'b01011_011111_01010;
        tomato_soup_dim[28][8] = 16'b01011_011111_01010;
        tomato_soup_dim[28][9] = 16'b01011_011111_01010;
        tomato_soup_dim[28][10] = 16'b01011_011111_01010;
        tomato_soup_dim[28][11] = 16'b01011_011111_01010;
        tomato_soup_dim[28][12] = 16'b01011_011111_01010;
        tomato_soup_dim[28][13] = 16'b01011_011111_01010;
        tomato_soup_dim[28][14] = 16'b01011_011111_01010;
        tomato_soup_dim[28][15] = 16'b01011_011111_01010;
        tomato_soup_dim[28][16] = 16'b01011_011111_01010;
        tomato_soup_dim[28][17] = 16'b01011_011111_01010;
        tomato_soup_dim[28][18] = 16'b01011_011111_01010;
        tomato_soup_dim[28][19] = 16'b01011_011111_01010;
        tomato_soup_dim[28][20] = 16'b01011_011111_01010;
        tomato_soup_dim[28][21] = 16'b01011_011111_01010;
        tomato_soup_dim[28][22] = 16'b01011_011111_01010;
        tomato_soup_dim[28][23] = 16'b01011_011111_01010;
        tomato_soup_dim[28][24] = 16'b01011_011111_01010;
        tomato_soup_dim[28][25] = 16'b01011_011111_01010;
        tomato_soup_dim[28][26] = 16'b01011_011111_01010;
        tomato_soup_dim[28][27] = 16'b01011_011111_01010;
        tomato_soup_dim[28][28] = 16'b01011_011111_01010;
        tomato_soup_dim[28][29] = 16'b01011_011111_01010;
        tomato_soup_dim[28][30] = 16'b01011_011111_01010;
        tomato_soup_dim[28][31] = 16'b01011_011111_01010;
        tomato_soup_dim[29][0] = 16'b01011_011111_01010;
        tomato_soup_dim[29][1] = 16'b01011_011111_01010;
        tomato_soup_dim[29][2] = 16'b01011_011111_01010;
        tomato_soup_dim[29][3] = 16'b01011_011111_01010;
        tomato_soup_dim[29][4] = 16'b01011_011111_01010;
        tomato_soup_dim[29][5] = 16'b01011_011111_01010;
        tomato_soup_dim[29][6] = 16'b01011_011111_01010;
        tomato_soup_dim[29][7] = 16'b01011_011111_01010;
        tomato_soup_dim[29][8] = 16'b01011_011111_01010;
        tomato_soup_dim[29][9] = 16'b01011_011111_01010;
        tomato_soup_dim[29][10] = 16'b01011_011111_01010;
        tomato_soup_dim[29][11] = 16'b01011_011111_01010;
        tomato_soup_dim[29][12] = 16'b01011_011111_01010;
        tomato_soup_dim[29][13] = 16'b01011_011111_01010;
        tomato_soup_dim[29][14] = 16'b01011_011111_01010;
        tomato_soup_dim[29][15] = 16'b01011_011111_01010;
        tomato_soup_dim[29][16] = 16'b01011_011111_01010;
        tomato_soup_dim[29][17] = 16'b01011_011111_01010;
        tomato_soup_dim[29][18] = 16'b01011_011111_01010;
        tomato_soup_dim[29][19] = 16'b01011_011111_01010;
        tomato_soup_dim[29][20] = 16'b01011_011111_01010;
        tomato_soup_dim[29][21] = 16'b01011_011111_01010;
        tomato_soup_dim[29][22] = 16'b01011_011111_01010;
        tomato_soup_dim[29][23] = 16'b01011_011111_01010;
        tomato_soup_dim[29][24] = 16'b01011_011111_01010;
        tomato_soup_dim[29][25] = 16'b01011_011111_01010;
        tomato_soup_dim[29][26] = 16'b01011_011111_01010;
        tomato_soup_dim[29][27] = 16'b01011_011111_01010;
        tomato_soup_dim[29][28] = 16'b01011_011111_01010;
        tomato_soup_dim[29][29] = 16'b01011_011111_01010;
        tomato_soup_dim[29][30] = 16'b01011_011111_01010;
        tomato_soup_dim[29][31] = 16'b01011_011111_01010;
        tomato_soup_dim[30][0] = 16'b01011_011111_01010;
        tomato_soup_dim[30][1] = 16'b01011_011111_01010;
        tomato_soup_dim[30][2] = 16'b01011_011111_01010;
        tomato_soup_dim[30][3] = 16'b01011_011111_01010;
        tomato_soup_dim[30][4] = 16'b01011_011111_01010;
        tomato_soup_dim[30][5] = 16'b01011_011111_01010;
        tomato_soup_dim[30][6] = 16'b01011_011111_01010;
        tomato_soup_dim[30][7] = 16'b01011_011111_01010;
        tomato_soup_dim[30][8] = 16'b01011_011111_01010;
        tomato_soup_dim[30][9] = 16'b01011_011111_01010;
        tomato_soup_dim[30][10] = 16'b01011_011111_01010;
        tomato_soup_dim[30][11] = 16'b01011_011111_01010;
        tomato_soup_dim[30][12] = 16'b01011_011111_01010;
        tomato_soup_dim[30][13] = 16'b01011_011111_01010;
        tomato_soup_dim[30][14] = 16'b01011_011111_01010;
        tomato_soup_dim[30][15] = 16'b01011_011111_01010;
        tomato_soup_dim[30][16] = 16'b01011_011111_01010;
        tomato_soup_dim[30][17] = 16'b01011_011111_01010;
        tomato_soup_dim[30][18] = 16'b01011_011111_01010;
        tomato_soup_dim[30][19] = 16'b01011_011111_01010;
        tomato_soup_dim[30][20] = 16'b01011_011111_01010;
        tomato_soup_dim[30][21] = 16'b01011_011111_01010;
        tomato_soup_dim[30][22] = 16'b01011_011111_01010;
        tomato_soup_dim[30][23] = 16'b01011_011111_01010;
        tomato_soup_dim[30][24] = 16'b01011_011111_01010;
        tomato_soup_dim[30][25] = 16'b01011_011111_01010;
        tomato_soup_dim[30][26] = 16'b01011_011111_01010;
        tomato_soup_dim[30][27] = 16'b01011_011111_01010;
        tomato_soup_dim[30][28] = 16'b01011_011111_01010;
        tomato_soup_dim[30][29] = 16'b01011_011111_01010;
        tomato_soup_dim[30][30] = 16'b01011_011111_01010;
        tomato_soup_dim[30][31] = 16'b01011_011111_01010;
        tomato_soup_dim[31][0] = 16'b01011_011111_01010;
        tomato_soup_dim[31][1] = 16'b01011_011111_01010;
        tomato_soup_dim[31][2] = 16'b01011_011111_01010;
        tomato_soup_dim[31][3] = 16'b01011_011111_01010;
        tomato_soup_dim[31][4] = 16'b01011_011111_01010;
        tomato_soup_dim[31][5] = 16'b01011_011111_01010;
        tomato_soup_dim[31][6] = 16'b01011_011111_01010;
        tomato_soup_dim[31][7] = 16'b01011_011111_01010;
        tomato_soup_dim[31][8] = 16'b01011_011111_01010;
        tomato_soup_dim[31][9] = 16'b01011_011111_01010;
        tomato_soup_dim[31][10] = 16'b01011_011111_01010;
        tomato_soup_dim[31][11] = 16'b01011_011111_01010;
        tomato_soup_dim[31][12] = 16'b01011_011111_01010;
        tomato_soup_dim[31][13] = 16'b01011_011111_01010;
        tomato_soup_dim[31][14] = 16'b01011_011111_01010;
        tomato_soup_dim[31][15] = 16'b01011_011111_01010;
        tomato_soup_dim[31][16] = 16'b01011_011111_01010;
        tomato_soup_dim[31][17] = 16'b01011_011111_01010;
        tomato_soup_dim[31][18] = 16'b01011_011111_01010;
        tomato_soup_dim[31][19] = 16'b01011_011111_01010;
        tomato_soup_dim[31][20] = 16'b01011_011111_01010;
        tomato_soup_dim[31][21] = 16'b01011_011111_01010;
        tomato_soup_dim[31][22] = 16'b01011_011111_01010;
        tomato_soup_dim[31][23] = 16'b01011_011111_01010;
        tomato_soup_dim[31][24] = 16'b01011_011111_01010;
        tomato_soup_dim[31][25] = 16'b01011_011111_01010;
        tomato_soup_dim[31][26] = 16'b01011_011111_01010;
        tomato_soup_dim[31][27] = 16'b01011_011111_01010;
        tomato_soup_dim[31][28] = 16'b01011_011111_01010;
        tomato_soup_dim[31][29] = 16'b01011_011111_01010;
        tomato_soup_dim[31][30] = 16'b01011_011111_01010;
        tomato_soup_dim[31][31] = 16'b01011_011111_01010;
        
        
        
        tomato_rice_dim[0][0] = 16'b01111_011000_01111;
        tomato_rice_dim[0][1] = 16'b01111_011000_01111;
        tomato_rice_dim[0][2] = 16'b01111_011000_01111;
        tomato_rice_dim[0][3] = 16'b01111_011000_01111;
        tomato_rice_dim[0][4] = 16'b01111_011000_01111;
        tomato_rice_dim[0][5] = 16'b01111_011000_01111;
        tomato_rice_dim[0][6] = 16'b01111_011000_01111;
        tomato_rice_dim[0][7] = 16'b01111_011000_01111;
        tomato_rice_dim[0][8] = 16'b01111_011000_01111;
        tomato_rice_dim[0][9] = 16'b01111_011000_01111;
        tomato_rice_dim[0][10] = 16'b01111_011000_01111;
        tomato_rice_dim[0][11] = 16'b01111_011000_01111;
        tomato_rice_dim[0][12] = 16'b01111_011000_01111;
        tomato_rice_dim[0][13] = 16'b01111_011000_01111;
        tomato_rice_dim[0][14] = 16'b01111_011000_01111;
        tomato_rice_dim[0][15] = 16'b01111_011000_01111;
        tomato_rice_dim[0][16] = 16'b01111_011000_01111;
        tomato_rice_dim[0][17] = 16'b01111_011000_01111;
        tomato_rice_dim[0][18] = 16'b01111_011000_01111;
        tomato_rice_dim[0][19] = 16'b01111_011000_01111;
        tomato_rice_dim[0][20] = 16'b01111_011000_01111;
        tomato_rice_dim[0][21] = 16'b01111_011000_01111;
        tomato_rice_dim[0][22] = 16'b01111_011000_01111;
        tomato_rice_dim[0][23] = 16'b01111_011000_01111;
        tomato_rice_dim[0][24] = 16'b01111_011000_01111;
        tomato_rice_dim[0][25] = 16'b01111_011000_01111;
        tomato_rice_dim[0][26] = 16'b01111_011000_01111;
        tomato_rice_dim[0][27] = 16'b01111_011000_01111;
        tomato_rice_dim[0][28] = 16'b01111_011000_01111;
        tomato_rice_dim[0][29] = 16'b01111_011000_01111;
        tomato_rice_dim[0][30] = 16'b01111_011000_01111;
        tomato_rice_dim[0][31] = 16'b01111_011000_01111;
        tomato_rice_dim[1][0] = 16'b01111_011000_01111;
        tomato_rice_dim[1][1] = 16'b01111_011000_01111;
        tomato_rice_dim[1][2] = 16'b01111_011000_01111;
        tomato_rice_dim[1][3] = 16'b01111_011000_01111;
        tomato_rice_dim[1][4] = 16'b01111_011000_01111;
        tomato_rice_dim[1][5] = 16'b01111_011000_01111;
        tomato_rice_dim[1][6] = 16'b01111_011000_01111;
        tomato_rice_dim[1][7] = 16'b01111_011000_01111;
        tomato_rice_dim[1][8] = 16'b01111_011000_01111;
        tomato_rice_dim[1][9] = 16'b01111_011000_01111;
        tomato_rice_dim[1][10] = 16'b01111_011000_01111;
        tomato_rice_dim[1][11] = 16'b01111_011000_01111;
        tomato_rice_dim[1][12] = 16'b01111_011000_01111;
        tomato_rice_dim[1][13] = 16'b01111_011000_01111;
        tomato_rice_dim[1][14] = 16'b01111_011000_01111;
        tomato_rice_dim[1][15] = 16'b01111_011000_01111;
        tomato_rice_dim[1][16] = 16'b01111_011000_01111;
        tomato_rice_dim[1][17] = 16'b01111_011000_01111;
        tomato_rice_dim[1][18] = 16'b01111_011000_01111;
        tomato_rice_dim[1][19] = 16'b01111_011000_01111;
        tomato_rice_dim[1][20] = 16'b01111_011000_01111;
        tomato_rice_dim[1][21] = 16'b01111_011000_01111;
        tomato_rice_dim[1][22] = 16'b01111_011000_01111;
        tomato_rice_dim[1][23] = 16'b01111_011000_01111;
        tomato_rice_dim[1][24] = 16'b01111_011000_01111;
        tomato_rice_dim[1][25] = 16'b01111_011000_01111;
        tomato_rice_dim[1][26] = 16'b01111_011000_01111;
        tomato_rice_dim[1][27] = 16'b01111_011000_01111;
        tomato_rice_dim[1][28] = 16'b01111_011000_01111;
        tomato_rice_dim[1][29] = 16'b01111_011000_01111;
        tomato_rice_dim[1][30] = 16'b01111_011000_01111;
        tomato_rice_dim[1][31] = 16'b01111_011000_01111;
        tomato_rice_dim[2][0] = 16'b01111_011000_01111;
        tomato_rice_dim[2][1] = 16'b01111_011000_01111;
        tomato_rice_dim[2][2] = 16'b01111_011000_01111;
        tomato_rice_dim[2][3] = 16'b01111_011000_01111;
        tomato_rice_dim[2][4] = 16'b01111_011000_01111;
        tomato_rice_dim[2][5] = 16'b01111_011000_01111;
        tomato_rice_dim[2][6] = 16'b01111_011000_01111;
        tomato_rice_dim[2][7] = 16'b01111_011000_01111;
        tomato_rice_dim[2][8] = 16'b01111_011000_01111;
        tomato_rice_dim[2][9] = 16'b01111_011000_01111;
        tomato_rice_dim[2][10] = 16'b01111_011000_01111;
        tomato_rice_dim[2][11] = 16'b01111_011000_01111;
        tomato_rice_dim[2][12] = 16'b01111_011000_01111;
        tomato_rice_dim[2][13] = 16'b01111_011000_01111;
        tomato_rice_dim[2][14] = 16'b01111_011000_01111;
        tomato_rice_dim[2][15] = 16'b01111_011000_01111;
        tomato_rice_dim[2][16] = 16'b01111_011000_01111;
        tomato_rice_dim[2][17] = 16'b01111_011000_01111;
        tomato_rice_dim[2][18] = 16'b01111_011000_01111;
        tomato_rice_dim[2][19] = 16'b01111_011000_01111;
        tomato_rice_dim[2][20] = 16'b01111_011000_01111;
        tomato_rice_dim[2][21] = 16'b01111_011000_01111;
        tomato_rice_dim[2][22] = 16'b01111_011000_01111;
        tomato_rice_dim[2][23] = 16'b01111_011000_01111;
        tomato_rice_dim[2][24] = 16'b01111_011000_01111;
        tomato_rice_dim[2][25] = 16'b01111_011000_01111;
        tomato_rice_dim[2][26] = 16'b01111_011000_01111;
        tomato_rice_dim[2][27] = 16'b01111_011000_01111;
        tomato_rice_dim[2][28] = 16'b01111_011000_01111;
        tomato_rice_dim[2][29] = 16'b01111_011000_01111;
        tomato_rice_dim[2][30] = 16'b01111_011000_01111;
        tomato_rice_dim[2][31] = 16'b01111_011000_01111;
        tomato_rice_dim[3][0] = 16'b01111_011000_01111;
        tomato_rice_dim[3][1] = 16'b01111_011000_01111;
        tomato_rice_dim[3][2] = 16'b01111_011000_01111;
        tomato_rice_dim[3][3] = 16'b01111_011000_01111;
        tomato_rice_dim[3][4] = 16'b01111_011000_01111;
        tomato_rice_dim[3][5] = 16'b01111_011000_01111;
        tomato_rice_dim[3][6] = 16'b01111_011000_01111;
        tomato_rice_dim[3][7] = 16'b01111_011000_01111;
        tomato_rice_dim[3][8] = 16'b01111_011000_01111;
        tomato_rice_dim[3][9] = 16'b01111_011000_01111;
        tomato_rice_dim[3][10] = 16'b01111_011000_01111;
        tomato_rice_dim[3][11] = 16'b01111_011000_01111;
        tomato_rice_dim[3][12] = 16'b01111_011000_01111;
        tomato_rice_dim[3][13] = 16'b01111_011000_01111;
        tomato_rice_dim[3][14] = 16'b01111_011000_01111;
        tomato_rice_dim[3][15] = 16'b01111_011000_01111;
        tomato_rice_dim[3][16] = 16'b01111_011000_01111;
        tomato_rice_dim[3][17] = 16'b01111_011000_01111;
        tomato_rice_dim[3][18] = 16'b01111_011000_01111;
        tomato_rice_dim[3][19] = 16'b01111_011000_01111;
        tomato_rice_dim[3][20] = 16'b01111_011000_01111;
        tomato_rice_dim[3][21] = 16'b01111_011000_01111;
        tomato_rice_dim[3][22] = 16'b01111_011000_01111;
        tomato_rice_dim[3][23] = 16'b01111_011000_01111;
        tomato_rice_dim[3][24] = 16'b01111_011000_01111;
        tomato_rice_dim[3][25] = 16'b01111_011000_01111;
        tomato_rice_dim[3][26] = 16'b01111_011000_01111;
        tomato_rice_dim[3][27] = 16'b01111_011000_01111;
        tomato_rice_dim[3][28] = 16'b01111_011000_01111;
        tomato_rice_dim[3][29] = 16'b01111_011000_01111;
        tomato_rice_dim[3][30] = 16'b01111_011000_01111;
        tomato_rice_dim[3][31] = 16'b01111_011000_01111;
        tomato_rice_dim[4][0] = 16'b01111_011000_01111;
        tomato_rice_dim[4][1] = 16'b01111_011000_01111;
        tomato_rice_dim[4][2] = 16'b01111_011000_01111;
        tomato_rice_dim[4][3] = 16'b01111_011000_01111;
        tomato_rice_dim[4][4] = 16'b01111_011000_01111;
        tomato_rice_dim[4][5] = 16'b01111_011000_01111;
        tomato_rice_dim[4][6] = 16'b01111_011000_01111;
        tomato_rice_dim[4][7] = 16'b01111_011000_01111;
        tomato_rice_dim[4][8] = 16'b01111_011000_01111;
        tomato_rice_dim[4][9] = 16'b01111_011000_01111;
        tomato_rice_dim[4][10] = 16'b01111_011000_01111;
        tomato_rice_dim[4][11] = 16'b01111_011000_01111;
        tomato_rice_dim[4][12] = 16'b01111_011000_01111;
        tomato_rice_dim[4][13] = 16'b01111_011000_01111;
        tomato_rice_dim[4][14] = 16'b01111_011000_01111;
        tomato_rice_dim[4][15] = 16'b01111_011000_01111;
        tomato_rice_dim[4][16] = 16'b01111_011000_01111;
        tomato_rice_dim[4][17] = 16'b01111_011000_01111;
        tomato_rice_dim[4][18] = 16'b01111_011000_01111;
        tomato_rice_dim[4][19] = 16'b01111_011000_01111;
        tomato_rice_dim[4][20] = 16'b01111_011000_01111;
        tomato_rice_dim[4][21] = 16'b01111_011000_01111;
        tomato_rice_dim[4][22] = 16'b01111_011000_01111;
        tomato_rice_dim[4][23] = 16'b01111_011000_01111;
        tomato_rice_dim[4][24] = 16'b01111_011000_01111;
        tomato_rice_dim[4][25] = 16'b01111_011000_01111;
        tomato_rice_dim[4][26] = 16'b01111_011000_01111;
        tomato_rice_dim[4][27] = 16'b01111_011000_01111;
        tomato_rice_dim[4][28] = 16'b01111_011000_01111;
        tomato_rice_dim[4][29] = 16'b01111_011000_01111;
        tomato_rice_dim[4][30] = 16'b01111_011000_01111;
        tomato_rice_dim[4][31] = 16'b01111_011000_01111;
        tomato_rice_dim[5][0] = 16'b01111_011000_01111;
        tomato_rice_dim[5][1] = 16'b01111_011000_01111;
        tomato_rice_dim[5][2] = 16'b01111_011000_01111;
        tomato_rice_dim[5][3] = 16'b01111_011000_01111;
        tomato_rice_dim[5][4] = 16'b01111_011000_01111;
        tomato_rice_dim[5][5] = 16'b01111_011000_01111;
        tomato_rice_dim[5][6] = 16'b01111_011000_01111;
        tomato_rice_dim[5][7] = 16'b01111_011000_01111;
        tomato_rice_dim[5][8] = 16'b01111_011000_01111;
        tomato_rice_dim[5][9] = 16'b01111_011000_01111;
        tomato_rice_dim[5][10] = 16'b01100_010100_00110;
        tomato_rice_dim[5][11] = 16'b01100_010100_00110;
        tomato_rice_dim[5][12] = 16'b01100_010100_00110;
        tomato_rice_dim[5][13] = 16'b01100_010100_00110;
        tomato_rice_dim[5][14] = 16'b01100_010100_00110;
        tomato_rice_dim[5][15] = 16'b01101_010110_00111;
        tomato_rice_dim[5][16] = 16'b01101_010101_00111;
        tomato_rice_dim[5][17] = 16'b01101_010101_00110;
        tomato_rice_dim[5][18] = 16'b01101_010101_00110;
        tomato_rice_dim[5][19] = 16'b01100_010101_00110;
        tomato_rice_dim[5][20] = 16'b01100_010101_00110;
        tomato_rice_dim[5][21] = 16'b01100_010101_00110;
        tomato_rice_dim[5][22] = 16'b01111_011000_01111;
        tomato_rice_dim[5][23] = 16'b01111_011000_01111;
        tomato_rice_dim[5][24] = 16'b01111_011000_01111;
        tomato_rice_dim[5][25] = 16'b01111_011000_01111;
        tomato_rice_dim[5][26] = 16'b01111_011000_01111;
        tomato_rice_dim[5][27] = 16'b01111_011000_01111;
        tomato_rice_dim[5][28] = 16'b01111_011000_01111;
        tomato_rice_dim[5][29] = 16'b01111_011000_01111;
        tomato_rice_dim[5][30] = 16'b01111_011000_01111;
        tomato_rice_dim[5][31] = 16'b01111_011000_01111;
        tomato_rice_dim[6][0] = 16'b01111_011000_01111;
        tomato_rice_dim[6][1] = 16'b01111_011000_01111;
        tomato_rice_dim[6][2] = 16'b01111_011000_01111;
        tomato_rice_dim[6][3] = 16'b01111_011000_01111;
        tomato_rice_dim[6][4] = 16'b01111_011000_01111;
        tomato_rice_dim[6][5] = 16'b01111_011000_01111;
        tomato_rice_dim[6][6] = 16'b01111_011000_01111;
        tomato_rice_dim[6][7] = 16'b01100_010100_00110;
        tomato_rice_dim[6][8] = 16'b01100_010100_00110;
        tomato_rice_dim[6][9] = 16'b01101_010111_00111;
        tomato_rice_dim[6][10] = 16'b01101_011000_01000;
        tomato_rice_dim[6][11] = 16'b01101_011000_01000;
        tomato_rice_dim[6][12] = 16'b01101_010111_01000;
        tomato_rice_dim[6][13] = 16'b01110_011000_01000;
        tomato_rice_dim[6][14] = 16'b01101_010111_01000;
        tomato_rice_dim[6][15] = 16'b01101_010110_00111;
        tomato_rice_dim[6][16] = 16'b01101_010111_01000;
        tomato_rice_dim[6][17] = 16'b01101_010111_01000;
        tomato_rice_dim[6][18] = 16'b01101_010111_01000;
        tomato_rice_dim[6][19] = 16'b01101_010111_01000;
        tomato_rice_dim[6][20] = 16'b01101_010111_01000;
        tomato_rice_dim[6][21] = 16'b01101_010110_00111;
        tomato_rice_dim[6][22] = 16'b01101_010101_00110;
        tomato_rice_dim[6][23] = 16'b01101_010101_00111;
        tomato_rice_dim[6][24] = 16'b01100_010100_00110;
        tomato_rice_dim[6][25] = 16'b01111_011000_01111;
        tomato_rice_dim[6][26] = 16'b01111_011000_01111;
        tomato_rice_dim[6][27] = 16'b01111_011000_01111;
        tomato_rice_dim[6][28] = 16'b01111_011000_01111;
        tomato_rice_dim[6][29] = 16'b01111_011000_01111;
        tomato_rice_dim[6][30] = 16'b01111_011000_01111;
        tomato_rice_dim[6][31] = 16'b01111_011000_01111;
        tomato_rice_dim[7][0] = 16'b01111_011000_01111;
        tomato_rice_dim[7][1] = 16'b01111_011000_01111;
        tomato_rice_dim[7][2] = 16'b01111_011000_01111;
        tomato_rice_dim[7][3] = 16'b01111_011000_01111;
        tomato_rice_dim[7][4] = 16'b01111_011000_01111;
        tomato_rice_dim[7][5] = 16'b01100_010100_00110;
        tomato_rice_dim[7][6] = 16'b01100_010100_00110;
        tomato_rice_dim[7][7] = 16'b01101_010111_01000;
        tomato_rice_dim[7][8] = 16'b01101_010111_01000;
        tomato_rice_dim[7][9] = 16'b01101_010111_01000;
        tomato_rice_dim[7][10] = 16'b01101_010111_00111;
        tomato_rice_dim[7][11] = 16'b01101_011000_01000;
        tomato_rice_dim[7][12] = 16'b01101_010111_01000;
        tomato_rice_dim[7][13] = 16'b01101_010111_01000;
        tomato_rice_dim[7][14] = 16'b01101_010111_01000;
        tomato_rice_dim[7][15] = 16'b01101_010110_00111;
        tomato_rice_dim[7][16] = 16'b01101_010110_00111;
        tomato_rice_dim[7][17] = 16'b01101_010111_00111;
        tomato_rice_dim[7][18] = 16'b01101_010110_00111;
        tomato_rice_dim[7][19] = 16'b01101_010110_00111;
        tomato_rice_dim[7][20] = 16'b01101_010111_00111;
        tomato_rice_dim[7][21] = 16'b01101_010111_01000;
        tomato_rice_dim[7][22] = 16'b01101_010111_00111;
        tomato_rice_dim[7][23] = 16'b01101_010111_01000;
        tomato_rice_dim[7][24] = 16'b01101_010111_01000;
        tomato_rice_dim[7][25] = 16'b01100_010100_00110;
        tomato_rice_dim[7][26] = 16'b01100_010100_00110;
        tomato_rice_dim[7][27] = 16'b01111_011000_01111;
        tomato_rice_dim[7][28] = 16'b01111_011000_01111;
        tomato_rice_dim[7][29] = 16'b01111_011000_01111;
        tomato_rice_dim[7][30] = 16'b01111_011000_01111;
        tomato_rice_dim[7][31] = 16'b01111_011000_01111;
        tomato_rice_dim[8][0] = 16'b01111_011000_01111;
        tomato_rice_dim[8][1] = 16'b01111_011000_01111;
        tomato_rice_dim[8][2] = 16'b01111_011000_01111;
        tomato_rice_dim[8][3] = 16'b01111_011000_01111;
        tomato_rice_dim[8][4] = 16'b01100_010011_00101;
        tomato_rice_dim[8][5] = 16'b01101_010111_00111;
        tomato_rice_dim[8][6] = 16'b01101_011000_01000;
        tomato_rice_dim[8][7] = 16'b01110_011000_01000;
        tomato_rice_dim[8][8] = 16'b01101_010111_00111;
        tomato_rice_dim[8][9] = 16'b01101_010110_00111;
        tomato_rice_dim[8][10] = 16'b01101_011000_01000;
        tomato_rice_dim[8][11] = 16'b01101_010111_01000;
        tomato_rice_dim[8][12] = 16'b01101_010101_00111;
        tomato_rice_dim[8][13] = 16'b01100_010100_00110;
        tomato_rice_dim[8][14] = 16'b01101_010100_00110;
        tomato_rice_dim[8][15] = 16'b01101_010100_00110;
        tomato_rice_dim[8][16] = 16'b01100_010100_00110;
        tomato_rice_dim[8][17] = 16'b01100_010011_00101;
        tomato_rice_dim[8][18] = 16'b01100_010010_00101;
        tomato_rice_dim[8][19] = 16'b01101_010101_00111;
        tomato_rice_dim[8][20] = 16'b01101_010111_01000;
        tomato_rice_dim[8][21] = 16'b01101_010111_00111;
        tomato_rice_dim[8][22] = 16'b01101_010111_00111;
        tomato_rice_dim[8][23] = 16'b01101_010111_01000;
        tomato_rice_dim[8][24] = 16'b01101_011000_01000;
        tomato_rice_dim[8][25] = 16'b01110_011000_01000;
        tomato_rice_dim[8][26] = 16'b01101_010111_01000;
        tomato_rice_dim[8][27] = 16'b01100_010100_00110;
        tomato_rice_dim[8][28] = 16'b01111_011000_01111;
        tomato_rice_dim[8][29] = 16'b01111_011000_01111;
        tomato_rice_dim[8][30] = 16'b01111_011000_01111;
        tomato_rice_dim[8][31] = 16'b01111_011000_01111;
        tomato_rice_dim[9][0] = 16'b01111_011000_01111;
        tomato_rice_dim[9][1] = 16'b01111_011000_01111;
        tomato_rice_dim[9][2] = 16'b01111_011000_01111;
        tomato_rice_dim[9][3] = 16'b01100_010100_00110;
        tomato_rice_dim[9][4] = 16'b01101_010111_01000;
        tomato_rice_dim[9][5] = 16'b01101_010111_01000;
        tomato_rice_dim[9][6] = 16'b01101_010111_01000;
        tomato_rice_dim[9][7] = 16'b01101_011000_01000;
        tomato_rice_dim[9][8] = 16'b01101_010111_01000;
        tomato_rice_dim[9][9] = 16'b01101_010101_00110;
        tomato_rice_dim[9][10] = 16'b01101_010101_00110;
        tomato_rice_dim[9][11] = 16'b01101_010101_00110;
        tomato_rice_dim[9][12] = 16'b01100_010000_00100;
        tomato_rice_dim[9][13] = 16'b01100_001101_00010;
        tomato_rice_dim[9][14] = 16'b01100_001011_00010;
        tomato_rice_dim[9][15] = 16'b01100_000111_00000;
        tomato_rice_dim[9][16] = 16'b01100_000111_00000;
        tomato_rice_dim[9][17] = 16'b01100_001011_00001;
        tomato_rice_dim[9][18] = 16'b01100_001100_00010;
        tomato_rice_dim[9][19] = 16'b01100_010010_00101;
        tomato_rice_dim[9][20] = 16'b01100_010100_00110;
        tomato_rice_dim[9][21] = 16'b01101_010101_00110;
        tomato_rice_dim[9][22] = 16'b01101_010101_00110;
        tomato_rice_dim[9][23] = 16'b01101_010111_00111;
        tomato_rice_dim[9][24] = 16'b01101_010111_01000;
        tomato_rice_dim[9][25] = 16'b01101_010111_01000;
        tomato_rice_dim[9][26] = 16'b01101_010111_01000;
        tomato_rice_dim[9][27] = 16'b01110_011000_01000;
        tomato_rice_dim[9][28] = 16'b01100_010101_00110;
        tomato_rice_dim[9][29] = 16'b01111_011000_01111;
        tomato_rice_dim[9][30] = 16'b01111_011000_01111;
        tomato_rice_dim[9][31] = 16'b01111_011000_01111;
        tomato_rice_dim[10][0] = 16'b01111_011000_01111;
        tomato_rice_dim[10][1] = 16'b01111_011000_01111;
        tomato_rice_dim[10][2] = 16'b01111_011000_01111;
        tomato_rice_dim[10][3] = 16'b01101_010111_01000;
        tomato_rice_dim[10][4] = 16'b01101_010111_01000;
        tomato_rice_dim[10][5] = 16'b01101_010111_01000;
        tomato_rice_dim[10][6] = 16'b01101_010111_00111;
        tomato_rice_dim[10][7] = 16'b01101_010101_00110;
        tomato_rice_dim[10][8] = 16'b01101_010100_00110;
        tomato_rice_dim[10][9] = 16'b01101_010000_00100;
        tomato_rice_dim[10][10] = 16'b01101_001101_00011;
        tomato_rice_dim[10][11] = 16'b01100_001000_00001;
        tomato_rice_dim[10][12] = 16'b01100_001000_00000;
        tomato_rice_dim[10][13] = 16'b01101_001001_00001;
        tomato_rice_dim[10][14] = 16'b01100_001001_00001;
        tomato_rice_dim[10][15] = 16'b01100_001000_00000;
        tomato_rice_dim[10][16] = 16'b01100_001001_00001;
        tomato_rice_dim[10][17] = 16'b01100_001001_00001;
        tomato_rice_dim[10][18] = 16'b01101_001010_00001;
        tomato_rice_dim[10][19] = 16'b01101_001010_00001;
        tomato_rice_dim[10][20] = 16'b01100_001001_00001;
        tomato_rice_dim[10][21] = 16'b01100_001000_00000;
        tomato_rice_dim[10][22] = 16'b01101_001110_00011;
        tomato_rice_dim[10][23] = 16'b01101_010101_00110;
        tomato_rice_dim[10][24] = 16'b01100_010100_00110;
        tomato_rice_dim[10][25] = 16'b01101_010111_01000;
        tomato_rice_dim[10][26] = 16'b01110_011000_01000;
        tomato_rice_dim[10][27] = 16'b01101_010111_01000;
        tomato_rice_dim[10][28] = 16'b01101_010111_01000;
        tomato_rice_dim[10][29] = 16'b01111_011000_01111;
        tomato_rice_dim[10][30] = 16'b01111_011000_01111;
        tomato_rice_dim[10][31] = 16'b01111_011000_01111;
        tomato_rice_dim[11][0] = 16'b01111_011000_01111;
        tomato_rice_dim[11][1] = 16'b01111_011000_01111;
        tomato_rice_dim[11][2] = 16'b01101_010101_00111;
        tomato_rice_dim[11][3] = 16'b01101_010111_01000;
        tomato_rice_dim[11][4] = 16'b01110_011000_01000;
        tomato_rice_dim[11][5] = 16'b01101_011000_01000;
        tomato_rice_dim[11][6] = 16'b01101_010101_00110;
        tomato_rice_dim[11][7] = 16'b01101_001110_00011;
        tomato_rice_dim[11][8] = 16'b01100_001000_00000;
        tomato_rice_dim[11][9] = 16'b01100_001000_00000;
        tomato_rice_dim[11][10] = 16'b01100_000111_00000;
        tomato_rice_dim[11][11] = 16'b01101_001010_00001;
        tomato_rice_dim[11][12] = 16'b01101_001010_00001;
        tomato_rice_dim[11][13] = 16'b01100_001001_00001;
        tomato_rice_dim[11][14] = 16'b01101_001011_00001;
        tomato_rice_dim[11][15] = 16'b01101_001010_00001;
        tomato_rice_dim[11][16] = 16'b01101_001010_00001;
        tomato_rice_dim[11][17] = 16'b01100_001001_00001;
        tomato_rice_dim[11][18] = 16'b01100_001001_00001;
        tomato_rice_dim[11][19] = 16'b01100_001001_00001;
        tomato_rice_dim[11][20] = 16'b01101_001001_00001;
        tomato_rice_dim[11][21] = 16'b01100_001001_00000;
        tomato_rice_dim[11][22] = 16'b01100_001001_00001;
        tomato_rice_dim[11][23] = 16'b01100_001000_00001;
        tomato_rice_dim[11][24] = 16'b01100_001111_00011;
        tomato_rice_dim[11][25] = 16'b01101_010100_00110;
        tomato_rice_dim[11][26] = 16'b01101_010111_01000;
        tomato_rice_dim[11][27] = 16'b01101_010111_00111;
        tomato_rice_dim[11][28] = 16'b01101_010111_00111;
        tomato_rice_dim[11][29] = 16'b01101_010110_00111;
        tomato_rice_dim[11][30] = 16'b01111_011000_01111;
        tomato_rice_dim[11][31] = 16'b01111_011000_01111;
        tomato_rice_dim[12][0] = 16'b01111_011000_01111;
        tomato_rice_dim[12][1] = 16'b01111_011000_01111;
        tomato_rice_dim[12][2] = 16'b01101_011000_01000;
        tomato_rice_dim[12][3] = 16'b01101_010111_01000;
        tomato_rice_dim[12][4] = 16'b01101_010111_01000;
        tomato_rice_dim[12][5] = 16'b01101_010101_00110;
        tomato_rice_dim[12][6] = 16'b01100_001101_00010;
        tomato_rice_dim[12][7] = 16'b01100_001000_00000;
        tomato_rice_dim[12][8] = 16'b01100_001000_00000;
        tomato_rice_dim[12][9] = 16'b01101_001001_00001;
        tomato_rice_dim[12][10] = 16'b01101_001001_00001;
        tomato_rice_dim[12][11] = 16'b01100_000111_00000;
        tomato_rice_dim[12][12] = 16'b01101_001001_00001;
        tomato_rice_dim[12][13] = 16'b01101_001001_00001;
        tomato_rice_dim[12][14] = 16'b01100_001001_00001;
        tomato_rice_dim[12][15] = 16'b01101_001010_00001;
        tomato_rice_dim[12][16] = 16'b01101_001001_00001;
        tomato_rice_dim[12][17] = 16'b01101_001001_00001;
        tomato_rice_dim[12][18] = 16'b01101_001010_00001;
        tomato_rice_dim[12][19] = 16'b01101_001010_00001;
        tomato_rice_dim[12][20] = 16'b01100_001000_00000;
        tomato_rice_dim[12][21] = 16'b01100_001000_00001;
        tomato_rice_dim[12][22] = 16'b01100_001001_00001;
        tomato_rice_dim[12][23] = 16'b01101_001001_00001;
        tomato_rice_dim[12][24] = 16'b01100_001000_00000;
        tomato_rice_dim[12][25] = 16'b01100_001100_00010;
        tomato_rice_dim[12][26] = 16'b01101_010100_00110;
        tomato_rice_dim[12][27] = 16'b01101_010111_01000;
        tomato_rice_dim[12][28] = 16'b01101_010111_00111;
        tomato_rice_dim[12][29] = 16'b01101_010111_01000;
        tomato_rice_dim[12][30] = 16'b01111_011000_01111;
        tomato_rice_dim[12][31] = 16'b01111_011000_01111;
        tomato_rice_dim[13][0] = 16'b01111_011000_01111;
        tomato_rice_dim[13][1] = 16'b01111_011000_01111;
        tomato_rice_dim[13][2] = 16'b01101_010111_01000;
        tomato_rice_dim[13][3] = 16'b01101_011000_01000;
        tomato_rice_dim[13][4] = 16'b01110_011000_01000;
        tomato_rice_dim[13][5] = 16'b01100_010100_00110;
        tomato_rice_dim[13][6] = 16'b01100_000111_00000;
        tomato_rice_dim[13][7] = 16'b01101_001001_00001;
        tomato_rice_dim[13][8] = 16'b01101_001001_00001;
        tomato_rice_dim[13][9] = 16'b01100_001000_00000;
        tomato_rice_dim[13][10] = 16'b01101_001001_00001;
        tomato_rice_dim[13][11] = 16'b01101_001001_00001;
        tomato_rice_dim[13][12] = 16'b01100_001000_00000;
        tomato_rice_dim[13][13] = 16'b01101_001010_00001;
        tomato_rice_dim[13][14] = 16'b01101_001010_00001;
        tomato_rice_dim[13][15] = 16'b01101_001001_00001;
        tomato_rice_dim[13][16] = 16'b01101_001011_00001;
        tomato_rice_dim[13][17] = 16'b01101_001010_00001;
        tomato_rice_dim[13][18] = 16'b01101_001011_00001;
        tomato_rice_dim[13][19] = 16'b01101_001001_00001;
        tomato_rice_dim[13][20] = 16'b01101_001010_00001;
        tomato_rice_dim[13][21] = 16'b01101_001001_00001;
        tomato_rice_dim[13][22] = 16'b01101_001001_00001;
        tomato_rice_dim[13][23] = 16'b01101_001100_00010;
        tomato_rice_dim[13][24] = 16'b01101_001001_00001;
        tomato_rice_dim[13][25] = 16'b01100_001000_00001;
        tomato_rice_dim[13][26] = 16'b01100_010100_00110;
        tomato_rice_dim[13][27] = 16'b01110_011000_01000;
        tomato_rice_dim[13][28] = 16'b01101_010111_01000;
        tomato_rice_dim[13][29] = 16'b01101_011000_01000;
        tomato_rice_dim[13][30] = 16'b01111_011000_01111;
        tomato_rice_dim[13][31] = 16'b01111_011000_01111;
        tomato_rice_dim[14][0] = 16'b01111_011000_01111;
        tomato_rice_dim[14][1] = 16'b01111_011000_01111;
        tomato_rice_dim[14][2] = 16'b01101_010111_01000;
        tomato_rice_dim[14][3] = 16'b01101_010111_01000;
        tomato_rice_dim[14][4] = 16'b01101_010111_01000;
        tomato_rice_dim[14][5] = 16'b01100_010100_00110;
        tomato_rice_dim[14][6] = 16'b01100_001001_00001;
        tomato_rice_dim[14][7] = 16'b01100_001001_00001;
        tomato_rice_dim[14][8] = 16'b01100_001001_00001;
        tomato_rice_dim[14][9] = 16'b01101_001001_00001;
        tomato_rice_dim[14][10] = 16'b01101_001001_00001;
        tomato_rice_dim[14][11] = 16'b01101_001011_00001;
        tomato_rice_dim[14][12] = 16'b01101_001010_00001;
        tomato_rice_dim[14][13] = 16'b01101_001010_00001;
        tomato_rice_dim[14][14] = 16'b01101_001100_00001;
        tomato_rice_dim[14][15] = 16'b01101_001010_00001;
        tomato_rice_dim[14][16] = 16'b01101_001010_00001;
        tomato_rice_dim[14][17] = 16'b01101_001010_00001;
        tomato_rice_dim[14][18] = 16'b01101_001001_00001;
        tomato_rice_dim[14][19] = 16'b01101_001010_00001;
        tomato_rice_dim[14][20] = 16'b01101_001010_00001;
        tomato_rice_dim[14][21] = 16'b01101_001011_00001;
        tomato_rice_dim[14][22] = 16'b01101_001010_00001;
        tomato_rice_dim[14][23] = 16'b01101_001001_00001;
        tomato_rice_dim[14][24] = 16'b01101_001001_00001;
        tomato_rice_dim[14][25] = 16'b01101_001010_00001;
        tomato_rice_dim[14][26] = 16'b01101_010101_00110;
        tomato_rice_dim[14][27] = 16'b01101_010111_01000;
        tomato_rice_dim[14][28] = 16'b01101_010110_00111;
        tomato_rice_dim[14][29] = 16'b01110_011000_01000;
        tomato_rice_dim[14][30] = 16'b01111_011000_01111;
        tomato_rice_dim[14][31] = 16'b01111_011000_01111;
        tomato_rice_dim[15][0] = 16'b01111_011000_01111;
        tomato_rice_dim[15][1] = 16'b01111_011000_01111;
        tomato_rice_dim[15][2] = 16'b01101_010111_01000;
        tomato_rice_dim[15][3] = 16'b01101_010111_01000;
        tomato_rice_dim[15][4] = 16'b01101_010111_01000;
        tomato_rice_dim[15][5] = 16'b01101_010101_00111;
        tomato_rice_dim[15][6] = 16'b01101_001011_00001;
        tomato_rice_dim[15][7] = 16'b01100_001000_00000;
        tomato_rice_dim[15][8] = 16'b01101_001001_00001;
        tomato_rice_dim[15][9] = 16'b01110_001100_00010;
        tomato_rice_dim[15][10] = 16'b01101_001100_00010;
        tomato_rice_dim[15][11] = 16'b01101_001001_00001;
        tomato_rice_dim[15][12] = 16'b01101_001100_00001;
        tomato_rice_dim[15][13] = 16'b01101_001010_00001;
        tomato_rice_dim[15][14] = 16'b01101_001011_00001;
        tomato_rice_dim[15][15] = 16'b01101_001010_00001;
        tomato_rice_dim[15][16] = 16'b01110_001101_00010;
        tomato_rice_dim[15][17] = 16'b01110_001101_00010;
        tomato_rice_dim[15][18] = 16'b01110_001100_00010;
        tomato_rice_dim[15][19] = 16'b01101_001011_00001;
        tomato_rice_dim[15][20] = 16'b01101_001001_00001;
        tomato_rice_dim[15][21] = 16'b01101_001010_00001;
        tomato_rice_dim[15][22] = 16'b01101_001011_00001;
        tomato_rice_dim[15][23] = 16'b01101_001100_00010;
        tomato_rice_dim[15][24] = 16'b01101_001001_00001;
        tomato_rice_dim[15][25] = 16'b01101_001010_00001;
        tomato_rice_dim[15][26] = 16'b01101_010111_00111;
        tomato_rice_dim[15][27] = 16'b01101_010111_00111;
        tomato_rice_dim[15][28] = 16'b01101_010110_00111;
        tomato_rice_dim[15][29] = 16'b01101_010111_01000;
        tomato_rice_dim[15][30] = 16'b01111_011000_01111;
        tomato_rice_dim[15][31] = 16'b01111_011000_01111;
        tomato_rice_dim[16][0] = 16'b01111_011000_01111;
        tomato_rice_dim[16][1] = 16'b01111_011000_01111;
        tomato_rice_dim[16][2] = 16'b01111_011000_01111;
        tomato_rice_dim[16][3] = 16'b01101_010110_00111;
        tomato_rice_dim[16][4] = 16'b01101_010111_00111;
        tomato_rice_dim[16][5] = 16'b01101_010110_00111;
        tomato_rice_dim[16][6] = 16'b01101_010001_00100;
        tomato_rice_dim[16][7] = 16'b01101_001010_00001;
        tomato_rice_dim[16][8] = 16'b01101_001010_00001;
        tomato_rice_dim[16][9] = 16'b01101_001010_00001;
        tomato_rice_dim[16][10] = 16'b01110_001100_00010;
        tomato_rice_dim[16][11] = 16'b01101_001011_00001;
        tomato_rice_dim[16][12] = 16'b01101_001100_00001;
        tomato_rice_dim[16][13] = 16'b01101_001100_00010;
        tomato_rice_dim[16][14] = 16'b01101_001011_00001;
        tomato_rice_dim[16][15] = 16'b01101_001011_00001;
        tomato_rice_dim[16][16] = 16'b01101_001010_00001;
        tomato_rice_dim[16][17] = 16'b01101_001100_00010;
        tomato_rice_dim[16][18] = 16'b01101_001010_00001;
        tomato_rice_dim[16][19] = 16'b01101_001011_00001;
        tomato_rice_dim[16][20] = 16'b01101_001010_00001;
        tomato_rice_dim[16][21] = 16'b01101_001001_00001;
        tomato_rice_dim[16][22] = 16'b01101_001010_00001;
        tomato_rice_dim[16][23] = 16'b01101_001011_00001;
        tomato_rice_dim[16][24] = 16'b01101_001010_00001;
        tomato_rice_dim[16][25] = 16'b01101_010000_00100;
        tomato_rice_dim[16][26] = 16'b01110_011000_01000;
        tomato_rice_dim[16][27] = 16'b01101_010111_00111;
        tomato_rice_dim[16][28] = 16'b01101_010111_01000;
        tomato_rice_dim[16][29] = 16'b01111_011000_01111;
        tomato_rice_dim[16][30] = 16'b01111_011000_01111;
        tomato_rice_dim[16][31] = 16'b01111_011000_01111;
        tomato_rice_dim[17][0] = 16'b01111_011000_01111;
        tomato_rice_dim[17][1] = 16'b01111_011000_01111;
        tomato_rice_dim[17][2] = 16'b01111_011000_01111;
        tomato_rice_dim[17][3] = 16'b01111_011000_01111;
        tomato_rice_dim[17][4] = 16'b01101_010110_00111;
        tomato_rice_dim[17][5] = 16'b01101_010110_00111;
        tomato_rice_dim[17][6] = 16'b01101_010111_00111;
        tomato_rice_dim[17][7] = 16'b01100_001000_00001;
        tomato_rice_dim[17][8] = 16'b01101_001010_00001;
        tomato_rice_dim[17][9] = 16'b01101_001011_00001;
        tomato_rice_dim[17][10] = 16'b01110_001100_00010;
        tomato_rice_dim[17][11] = 16'b01101_001011_00001;
        tomato_rice_dim[17][12] = 16'b01101_001010_00001;
        tomato_rice_dim[17][13] = 16'b01101_001100_00010;
        tomato_rice_dim[17][14] = 16'b01110_001111_00011;
        tomato_rice_dim[17][15] = 16'b01101_001100_00010;
        tomato_rice_dim[17][16] = 16'b01101_001011_00001;
        tomato_rice_dim[17][17] = 16'b01101_001011_00001;
        tomato_rice_dim[17][18] = 16'b01101_001100_00010;
        tomato_rice_dim[17][19] = 16'b01101_001011_00001;
        tomato_rice_dim[17][20] = 16'b01101_001011_00001;
        tomato_rice_dim[17][21] = 16'b01101_001100_00010;
        tomato_rice_dim[17][22] = 16'b01101_001011_00001;
        tomato_rice_dim[17][23] = 16'b01100_001000_00000;
        tomato_rice_dim[17][24] = 16'b01101_001010_00001;
        tomato_rice_dim[17][25] = 16'b01101_010110_00111;
        tomato_rice_dim[17][26] = 16'b01101_010111_00111;
        tomato_rice_dim[17][27] = 16'b01101_011000_01000;
        tomato_rice_dim[17][28] = 16'b01111_011000_01111;
        tomato_rice_dim[17][29] = 16'b01111_011000_01111;
        tomato_rice_dim[17][30] = 16'b01111_011000_01111;
        tomato_rice_dim[17][31] = 16'b01111_011000_01111;
        tomato_rice_dim[18][0] = 16'b01111_011000_01111;
        tomato_rice_dim[18][1] = 16'b01111_011000_01111;
        tomato_rice_dim[18][2] = 16'b01111_011000_01111;
        tomato_rice_dim[18][3] = 16'b01111_011000_01111;
        tomato_rice_dim[18][4] = 16'b01111_011000_01111;
        tomato_rice_dim[18][5] = 16'b01101_010110_00111;
        tomato_rice_dim[18][6] = 16'b01101_010110_00111;
        tomato_rice_dim[18][7] = 16'b01101_001010_00001;
        tomato_rice_dim[18][8] = 16'b01101_001001_00001;
        tomato_rice_dim[18][9] = 16'b01101_001011_00001;
        tomato_rice_dim[18][10] = 16'b01101_001001_00001;
        tomato_rice_dim[18][11] = 16'b01101_001011_00001;
        tomato_rice_dim[18][12] = 16'b01101_001100_00010;
        tomato_rice_dim[18][13] = 16'b01101_001101_00010;
        tomato_rice_dim[18][14] = 16'b01101_001100_00010;
        tomato_rice_dim[18][15] = 16'b01101_001011_00001;
        tomato_rice_dim[18][16] = 16'b01110_001101_00010;
        tomato_rice_dim[18][17] = 16'b01101_001011_00001;
        tomato_rice_dim[18][18] = 16'b01101_001100_00010;
        tomato_rice_dim[18][19] = 16'b01110_001101_00010;
        tomato_rice_dim[18][20] = 16'b01101_001011_00001;
        tomato_rice_dim[18][21] = 16'b01101_001001_00001;
        tomato_rice_dim[18][22] = 16'b01101_001010_00001;
        tomato_rice_dim[18][23] = 16'b01101_001011_00001;
        tomato_rice_dim[18][24] = 16'b01101_001010_00001;
        tomato_rice_dim[18][25] = 16'b01101_010110_00111;
        tomato_rice_dim[18][26] = 16'b01101_010111_00111;
        tomato_rice_dim[18][27] = 16'b01111_011000_01111;
        tomato_rice_dim[18][28] = 16'b01111_011000_01111;
        tomato_rice_dim[18][29] = 16'b01111_011000_01111;
        tomato_rice_dim[18][30] = 16'b01111_011000_01111;
        tomato_rice_dim[18][31] = 16'b01111_011000_01111;
        tomato_rice_dim[19][0] = 16'b01111_011000_01111;
        tomato_rice_dim[19][1] = 16'b01111_011000_01111;
        tomato_rice_dim[19][2] = 16'b01111_011000_01111;
        tomato_rice_dim[19][3] = 16'b01111_011000_01111;
        tomato_rice_dim[19][4] = 16'b01111_011000_01111;
        tomato_rice_dim[19][5] = 16'b01111_011000_01111;
        tomato_rice_dim[19][6] = 16'b01111_011000_01111;
        tomato_rice_dim[19][7] = 16'b01110_010010_00101;
        tomato_rice_dim[19][8] = 16'b01101_001010_00001;
        tomato_rice_dim[19][9] = 16'b01101_001011_00001;
        tomato_rice_dim[19][10] = 16'b01101_001100_00001;
        tomato_rice_dim[19][11] = 16'b01101_001100_00010;
        tomato_rice_dim[19][12] = 16'b01101_001010_00001;
        tomato_rice_dim[19][13] = 16'b01101_001100_00010;
        tomato_rice_dim[19][14] = 16'b01110_001111_00011;
        tomato_rice_dim[19][15] = 16'b01101_001100_00010;
        tomato_rice_dim[19][16] = 16'b01101_001100_00010;
        tomato_rice_dim[19][17] = 16'b01101_001100_00010;
        tomato_rice_dim[19][18] = 16'b01101_001100_00010;
        tomato_rice_dim[19][19] = 16'b01101_001011_00001;
        tomato_rice_dim[19][20] = 16'b01101_001100_00001;
        tomato_rice_dim[19][21] = 16'b01101_001001_00001;
        tomato_rice_dim[19][22] = 16'b01101_001010_00001;
        tomato_rice_dim[19][23] = 16'b01101_001011_00001;
        tomato_rice_dim[19][24] = 16'b01110_010010_00100;
        tomato_rice_dim[19][25] = 16'b01111_011000_01111;
        tomato_rice_dim[19][26] = 16'b01111_011000_01111;
        tomato_rice_dim[19][27] = 16'b01111_011000_01111;
        tomato_rice_dim[19][28] = 16'b01111_011000_01111;
        tomato_rice_dim[19][29] = 16'b01111_011000_01111;
        tomato_rice_dim[19][30] = 16'b01111_011000_01111;
        tomato_rice_dim[19][31] = 16'b01111_011000_01111;
        tomato_rice_dim[20][0] = 16'b01111_011000_01111;
        tomato_rice_dim[20][1] = 16'b01111_011000_01111;
        tomato_rice_dim[20][2] = 16'b01111_011000_01111;
        tomato_rice_dim[20][3] = 16'b01111_011000_01111;
        tomato_rice_dim[20][4] = 16'b01111_011000_01111;
        tomato_rice_dim[20][5] = 16'b01111_011000_01111;
        tomato_rice_dim[20][6] = 16'b01111_011000_01111;
        tomato_rice_dim[20][7] = 16'b01111_011000_01111;
        tomato_rice_dim[20][8] = 16'b01101_001100_00010;
        tomato_rice_dim[20][9] = 16'b01101_001010_00001;
        tomato_rice_dim[20][10] = 16'b01101_001011_00001;
        tomato_rice_dim[20][11] = 16'b01101_001100_00001;
        tomato_rice_dim[20][12] = 16'b01101_001100_00010;
        tomato_rice_dim[20][13] = 16'b01101_001100_00010;
        tomato_rice_dim[20][14] = 16'b01101_001011_00001;
        tomato_rice_dim[20][15] = 16'b01101_001100_00001;
        tomato_rice_dim[20][16] = 16'b01110_001110_00010;
        tomato_rice_dim[20][17] = 16'b01101_001100_00010;
        tomato_rice_dim[20][18] = 16'b01101_001011_00001;
        tomato_rice_dim[20][19] = 16'b01110_001110_00010;
        tomato_rice_dim[20][20] = 16'b01101_001100_00010;
        tomato_rice_dim[20][21] = 16'b01101_001011_00001;
        tomato_rice_dim[20][22] = 16'b01101_001001_00001;
        tomato_rice_dim[20][23] = 16'b01101_001011_00001;
        tomato_rice_dim[20][24] = 16'b01111_011000_01111;
        tomato_rice_dim[20][25] = 16'b01111_011000_01111;
        tomato_rice_dim[20][26] = 16'b01111_011000_01111;
        tomato_rice_dim[20][27] = 16'b01111_011000_01111;
        tomato_rice_dim[20][28] = 16'b01111_011000_01111;
        tomato_rice_dim[20][29] = 16'b01111_011000_01111;
        tomato_rice_dim[20][30] = 16'b01111_011000_01111;
        tomato_rice_dim[20][31] = 16'b01111_011000_01111;
        tomato_rice_dim[21][0] = 16'b01111_011000_01111;
        tomato_rice_dim[21][1] = 16'b01111_011000_01111;
        tomato_rice_dim[21][2] = 16'b01111_011000_01111;
        tomato_rice_dim[21][3] = 16'b01111_011000_01111;
        tomato_rice_dim[21][4] = 16'b01111_011000_01111;
        tomato_rice_dim[21][5] = 16'b01111_011000_01111;
        tomato_rice_dim[21][6] = 16'b01111_011000_01111;
        tomato_rice_dim[21][7] = 16'b01111_011000_01111;
        tomato_rice_dim[21][8] = 16'b01111_011000_01111;
        tomato_rice_dim[21][9] = 16'b01101_001100_00010;
        tomato_rice_dim[21][10] = 16'b01101_001011_00001;
        tomato_rice_dim[21][11] = 16'b01110_001101_00010;
        tomato_rice_dim[21][12] = 16'b01110_001101_00010;
        tomato_rice_dim[21][13] = 16'b01101_001010_00001;
        tomato_rice_dim[21][14] = 16'b01101_001100_00001;
        tomato_rice_dim[21][15] = 16'b01110_001110_00010;
        tomato_rice_dim[21][16] = 16'b01110_001110_00010;
        tomato_rice_dim[21][17] = 16'b01101_001011_00001;
        tomato_rice_dim[21][18] = 16'b01110_001101_00010;
        tomato_rice_dim[21][19] = 16'b01101_001011_00001;
        tomato_rice_dim[21][20] = 16'b01110_001100_00010;
        tomato_rice_dim[21][21] = 16'b01110_001101_00010;
        tomato_rice_dim[21][22] = 16'b01101_001011_00001;
        tomato_rice_dim[21][23] = 16'b01111_011000_01111;
        tomato_rice_dim[21][24] = 16'b01111_011000_01111;
        tomato_rice_dim[21][25] = 16'b01111_011000_01111;
        tomato_rice_dim[21][26] = 16'b01111_011000_01111;
        tomato_rice_dim[21][27] = 16'b01111_011000_01111;
        tomato_rice_dim[21][28] = 16'b01111_011000_01111;
        tomato_rice_dim[21][29] = 16'b01111_011000_01111;
        tomato_rice_dim[21][30] = 16'b01111_011000_01111;
        tomato_rice_dim[21][31] = 16'b01111_011000_01111;
        tomato_rice_dim[22][0] = 16'b01111_011000_01111;
        tomato_rice_dim[22][1] = 16'b01111_011000_01111;
        tomato_rice_dim[22][2] = 16'b01111_011000_01111;
        tomato_rice_dim[22][3] = 16'b01111_011000_01111;
        tomato_rice_dim[22][4] = 16'b01111_011000_01111;
        tomato_rice_dim[22][5] = 16'b01111_011000_01111;
        tomato_rice_dim[22][6] = 16'b01111_011000_01111;
        tomato_rice_dim[22][7] = 16'b01111_011000_01111;
        tomato_rice_dim[22][8] = 16'b01111_011000_01111;
        tomato_rice_dim[22][9] = 16'b01111_011000_01111;
        tomato_rice_dim[22][10] = 16'b01110_001011_00001;
        tomato_rice_dim[22][11] = 16'b01101_001011_00001;
        tomato_rice_dim[22][12] = 16'b01110_001101_00010;
        tomato_rice_dim[22][13] = 16'b01110_001101_00010;
        tomato_rice_dim[22][14] = 16'b01101_001011_00001;
        tomato_rice_dim[22][15] = 16'b01101_001100_00001;
        tomato_rice_dim[22][16] = 16'b01110_001100_00010;
        tomato_rice_dim[22][17] = 16'b01110_001100_00010;
        tomato_rice_dim[22][18] = 16'b01110_001110_00010;
        tomato_rice_dim[22][19] = 16'b01101_001100_00010;
        tomato_rice_dim[22][20] = 16'b01101_001001_00001;
        tomato_rice_dim[22][21] = 16'b01101_001010_00001;
        tomato_rice_dim[22][22] = 16'b01110_010000_00011;
        tomato_rice_dim[22][23] = 16'b01111_011000_01111;
        tomato_rice_dim[22][24] = 16'b01111_011000_01111;
        tomato_rice_dim[22][25] = 16'b01111_011000_01111;
        tomato_rice_dim[22][26] = 16'b01111_011000_01111;
        tomato_rice_dim[22][27] = 16'b01111_011000_01111;
        tomato_rice_dim[22][28] = 16'b01111_011000_01111;
        tomato_rice_dim[22][29] = 16'b01111_011000_01111;
        tomato_rice_dim[22][30] = 16'b01111_011000_01111;
        tomato_rice_dim[22][31] = 16'b01111_011000_01111;
        tomato_rice_dim[23][0] = 16'b01111_011000_01111;
        tomato_rice_dim[23][1] = 16'b01111_011000_01111;
        tomato_rice_dim[23][2] = 16'b01111_011000_01111;
        tomato_rice_dim[23][3] = 16'b01111_011000_01111;
        tomato_rice_dim[23][4] = 16'b01111_011000_01111;
        tomato_rice_dim[23][5] = 16'b01111_011000_01111;
        tomato_rice_dim[23][6] = 16'b01111_011000_01111;
        tomato_rice_dim[23][7] = 16'b01111_011000_01111;
        tomato_rice_dim[23][8] = 16'b01111_011000_01111;
        tomato_rice_dim[23][9] = 16'b01111_011000_01111;
        tomato_rice_dim[23][10] = 16'b01111_011000_01111;
        tomato_rice_dim[23][11] = 16'b01110_010000_00100;
        tomato_rice_dim[23][12] = 16'b01110_001101_00010;
        tomato_rice_dim[23][13] = 16'b01101_001011_00001;
        tomato_rice_dim[23][14] = 16'b01110_001100_00010;
        tomato_rice_dim[23][15] = 16'b01101_001011_00001;
        tomato_rice_dim[23][16] = 16'b01110_001100_00010;
        tomato_rice_dim[23][17] = 16'b01110_001100_00010;
        tomato_rice_dim[23][18] = 16'b01110_001100_00010;
        tomato_rice_dim[23][19] = 16'b01101_001011_00001;
        tomato_rice_dim[23][20] = 16'b01101_001011_00001;
        tomato_rice_dim[23][21] = 16'b01111_011000_01111;
        tomato_rice_dim[23][22] = 16'b01111_011000_01111;
        tomato_rice_dim[23][23] = 16'b01111_011000_01111;
        tomato_rice_dim[23][24] = 16'b01111_011000_01111;
        tomato_rice_dim[23][25] = 16'b01111_011000_01111;
        tomato_rice_dim[23][26] = 16'b01111_011000_01111;
        tomato_rice_dim[23][27] = 16'b01111_011000_01111;
        tomato_rice_dim[23][28] = 16'b01111_011000_01111;
        tomato_rice_dim[23][29] = 16'b01111_011000_01111;
        tomato_rice_dim[23][30] = 16'b01111_011000_01111;
        tomato_rice_dim[23][31] = 16'b01111_011000_01111;
        tomato_rice_dim[24][0] = 16'b01111_011000_01111;
        tomato_rice_dim[24][1] = 16'b01111_011000_01111;
        tomato_rice_dim[24][2] = 16'b01111_011000_01111;
        tomato_rice_dim[24][3] = 16'b01111_011000_01111;
        tomato_rice_dim[24][4] = 16'b01111_011000_01111;
        tomato_rice_dim[24][5] = 16'b01111_011000_01111;
        tomato_rice_dim[24][6] = 16'b01111_011000_01111;
        tomato_rice_dim[24][7] = 16'b01111_011000_01111;
        tomato_rice_dim[24][8] = 16'b01111_011000_01111;
        tomato_rice_dim[24][9] = 16'b01111_011000_01111;
        tomato_rice_dim[24][10] = 16'b01111_011000_01111;
        tomato_rice_dim[24][11] = 16'b01111_011000_01111;
        tomato_rice_dim[24][12] = 16'b01111_011000_01111;
        tomato_rice_dim[24][13] = 16'b01110_001101_00010;
        tomato_rice_dim[24][14] = 16'b01101_001010_00001;
        tomato_rice_dim[24][15] = 16'b01110_001101_00010;
        tomato_rice_dim[24][16] = 16'b01101_001010_00001;
        tomato_rice_dim[24][17] = 16'b01110_001101_00010;
        tomato_rice_dim[24][18] = 16'b01101_001010_00001;
        tomato_rice_dim[24][19] = 16'b01111_011000_01111;
        tomato_rice_dim[24][20] = 16'b01111_011000_01111;
        tomato_rice_dim[24][21] = 16'b01111_011000_01111;
        tomato_rice_dim[24][22] = 16'b01111_011000_01111;
        tomato_rice_dim[24][23] = 16'b01111_011000_01111;
        tomato_rice_dim[24][24] = 16'b01111_011000_01111;
        tomato_rice_dim[24][25] = 16'b01111_011000_01111;
        tomato_rice_dim[24][26] = 16'b01111_011000_01111;
        tomato_rice_dim[24][27] = 16'b01111_011000_01111;
        tomato_rice_dim[24][28] = 16'b01111_011000_01111;
        tomato_rice_dim[24][29] = 16'b01111_011000_01111;
        tomato_rice_dim[24][30] = 16'b01111_011000_01111;
        tomato_rice_dim[24][31] = 16'b01111_011000_01111;
        tomato_rice_dim[25][0] = 16'b01111_011000_01111;
        tomato_rice_dim[25][1] = 16'b01111_011000_01111;
        tomato_rice_dim[25][2] = 16'b01111_011000_01111;
        tomato_rice_dim[25][3] = 16'b01111_011000_01111;
        tomato_rice_dim[25][4] = 16'b01111_011000_01111;
        tomato_rice_dim[25][5] = 16'b01111_011000_01111;
        tomato_rice_dim[25][6] = 16'b01111_011000_01111;
        tomato_rice_dim[25][7] = 16'b01111_011000_01111;
        tomato_rice_dim[25][8] = 16'b01111_011000_01111;
        tomato_rice_dim[25][9] = 16'b01111_011000_01111;
        tomato_rice_dim[25][10] = 16'b01111_011000_01111;
        tomato_rice_dim[25][11] = 16'b01111_011000_01111;
        tomato_rice_dim[25][12] = 16'b01111_011000_01111;
        tomato_rice_dim[25][13] = 16'b01111_011000_01111;
        tomato_rice_dim[25][14] = 16'b01111_011000_01111;
        tomato_rice_dim[25][15] = 16'b01111_011000_01111;
        tomato_rice_dim[25][16] = 16'b01111_011000_01111;
        tomato_rice_dim[25][17] = 16'b01111_011000_01111;
        tomato_rice_dim[25][18] = 16'b01111_011000_01111;
        tomato_rice_dim[25][19] = 16'b01111_011000_01111;
        tomato_rice_dim[25][20] = 16'b01111_011000_01111;
        tomato_rice_dim[25][21] = 16'b01111_011000_01111;
        tomato_rice_dim[25][22] = 16'b01111_011000_01111;
        tomato_rice_dim[25][23] = 16'b01111_011000_01111;
        tomato_rice_dim[25][24] = 16'b01111_011000_01111;
        tomato_rice_dim[25][25] = 16'b01111_011000_01111;
        tomato_rice_dim[25][26] = 16'b01111_011000_01111;
        tomato_rice_dim[25][27] = 16'b01111_011000_01111;
        tomato_rice_dim[25][28] = 16'b01111_011000_01111;
        tomato_rice_dim[25][29] = 16'b01111_011000_01111;
        tomato_rice_dim[25][30] = 16'b01111_011000_01111;
        tomato_rice_dim[25][31] = 16'b01111_011000_01111;
        tomato_rice_dim[26][0] = 16'b01111_011000_01111;
        tomato_rice_dim[26][1] = 16'b01111_011000_01111;
        tomato_rice_dim[26][2] = 16'b01111_011000_01111;
        tomato_rice_dim[26][3] = 16'b01111_011000_01111;
        tomato_rice_dim[26][4] = 16'b01111_011000_01111;
        tomato_rice_dim[26][5] = 16'b01111_011000_01111;
        tomato_rice_dim[26][6] = 16'b01111_011000_01111;
        tomato_rice_dim[26][7] = 16'b01111_011000_01111;
        tomato_rice_dim[26][8] = 16'b01111_011000_01111;
        tomato_rice_dim[26][9] = 16'b01111_011000_01111;
        tomato_rice_dim[26][10] = 16'b01111_011000_01111;
        tomato_rice_dim[26][11] = 16'b01111_011000_01111;
        tomato_rice_dim[26][12] = 16'b01111_011000_01111;
        tomato_rice_dim[26][13] = 16'b01111_011000_01111;
        tomato_rice_dim[26][14] = 16'b01111_011000_01111;
        tomato_rice_dim[26][15] = 16'b01111_011000_01111;
        tomato_rice_dim[26][16] = 16'b01111_011000_01111;
        tomato_rice_dim[26][17] = 16'b01111_011000_01111;
        tomato_rice_dim[26][18] = 16'b01111_011000_01111;
        tomato_rice_dim[26][19] = 16'b01111_011000_01111;
        tomato_rice_dim[26][20] = 16'b01111_011000_01111;
        tomato_rice_dim[26][21] = 16'b01111_011000_01111;
        tomato_rice_dim[26][22] = 16'b01111_011000_01111;
        tomato_rice_dim[26][23] = 16'b01111_011000_01111;
        tomato_rice_dim[26][24] = 16'b01111_011000_01111;
        tomato_rice_dim[26][25] = 16'b01111_011000_01111;
        tomato_rice_dim[26][26] = 16'b01111_011000_01111;
        tomato_rice_dim[26][27] = 16'b01111_011000_01111;
        tomato_rice_dim[26][28] = 16'b01111_011000_01111;
        tomato_rice_dim[26][29] = 16'b01111_011000_01111;
        tomato_rice_dim[26][30] = 16'b01111_011000_01111;
        tomato_rice_dim[26][31] = 16'b01111_011000_01111;
        tomato_rice_dim[27][0] = 16'b01111_011000_01111;
        tomato_rice_dim[27][1] = 16'b01111_011000_01111;
        tomato_rice_dim[27][2] = 16'b01111_011000_01111;
        tomato_rice_dim[27][3] = 16'b01111_011000_01111;
        tomato_rice_dim[27][4] = 16'b01111_011000_01111;
        tomato_rice_dim[27][5] = 16'b01111_011000_01111;
        tomato_rice_dim[27][6] = 16'b01111_011000_01111;
        tomato_rice_dim[27][7] = 16'b01111_011000_01111;
        tomato_rice_dim[27][8] = 16'b01111_011000_01111;
        tomato_rice_dim[27][9] = 16'b01111_011000_01111;
        tomato_rice_dim[27][10] = 16'b01111_011000_01111;
        tomato_rice_dim[27][11] = 16'b01111_011000_01111;
        tomato_rice_dim[27][12] = 16'b01111_011000_01111;
        tomato_rice_dim[27][13] = 16'b01111_011000_01111;
        tomato_rice_dim[27][14] = 16'b01111_011000_01111;
        tomato_rice_dim[27][15] = 16'b01111_011000_01111;
        tomato_rice_dim[27][16] = 16'b01111_011000_01111;
        tomato_rice_dim[27][17] = 16'b01111_011000_01111;
        tomato_rice_dim[27][18] = 16'b01111_011000_01111;
        tomato_rice_dim[27][19] = 16'b01111_011000_01111;
        tomato_rice_dim[27][20] = 16'b01111_011000_01111;
        tomato_rice_dim[27][21] = 16'b01111_011000_01111;
        tomato_rice_dim[27][22] = 16'b01111_011000_01111;
        tomato_rice_dim[27][23] = 16'b01111_011000_01111;
        tomato_rice_dim[27][24] = 16'b01111_011000_01111;
        tomato_rice_dim[27][25] = 16'b01111_011000_01111;
        tomato_rice_dim[27][26] = 16'b01111_011000_01111;
        tomato_rice_dim[27][27] = 16'b01111_011000_01111;
        tomato_rice_dim[27][28] = 16'b01111_011000_01111;
        tomato_rice_dim[27][29] = 16'b01111_011000_01111;
        tomato_rice_dim[27][30] = 16'b01111_011000_01111;
        tomato_rice_dim[27][31] = 16'b01111_011000_01111;
        tomato_rice_dim[28][0] = 16'b01111_011000_01111;
        tomato_rice_dim[28][1] = 16'b01111_011000_01111;
        tomato_rice_dim[28][2] = 16'b01111_011000_01111;
        tomato_rice_dim[28][3] = 16'b01111_011000_01111;
        tomato_rice_dim[28][4] = 16'b01111_011000_01111;
        tomato_rice_dim[28][5] = 16'b01111_011000_01111;
        tomato_rice_dim[28][6] = 16'b01111_011000_01111;
        tomato_rice_dim[28][7] = 16'b01111_011000_01111;
        tomato_rice_dim[28][8] = 16'b01111_011000_01111;
        tomato_rice_dim[28][9] = 16'b01111_011000_01111;
        tomato_rice_dim[28][10] = 16'b01111_011000_01111;
        tomato_rice_dim[28][11] = 16'b01111_011000_01111;
        tomato_rice_dim[28][12] = 16'b01111_011000_01111;
        tomato_rice_dim[28][13] = 16'b01111_011000_01111;
        tomato_rice_dim[28][14] = 16'b01111_011000_01111;
        tomato_rice_dim[28][15] = 16'b01111_011000_01111;
        tomato_rice_dim[28][16] = 16'b01111_011000_01111;
        tomato_rice_dim[28][17] = 16'b01111_011000_01111;
        tomato_rice_dim[28][18] = 16'b01111_011000_01111;
        tomato_rice_dim[28][19] = 16'b01111_011000_01111;
        tomato_rice_dim[28][20] = 16'b01111_011000_01111;
        tomato_rice_dim[28][21] = 16'b01111_011000_01111;
        tomato_rice_dim[28][22] = 16'b01111_011000_01111;
        tomato_rice_dim[28][23] = 16'b01111_011000_01111;
        tomato_rice_dim[28][24] = 16'b01111_011000_01111;
        tomato_rice_dim[28][25] = 16'b01111_011000_01111;
        tomato_rice_dim[28][26] = 16'b01111_011000_01111;
        tomato_rice_dim[28][27] = 16'b01111_011000_01111;
        tomato_rice_dim[28][28] = 16'b01111_011000_01111;
        tomato_rice_dim[28][29] = 16'b01111_011000_01111;
        tomato_rice_dim[28][30] = 16'b01111_011000_01111;
        tomato_rice_dim[28][31] = 16'b01111_011000_01111;
        tomato_rice_dim[29][0] = 16'b01111_011000_01111;
        tomato_rice_dim[29][1] = 16'b01111_011000_01111;
        tomato_rice_dim[29][2] = 16'b01111_011000_01111;
        tomato_rice_dim[29][3] = 16'b01111_011000_01111;
        tomato_rice_dim[29][4] = 16'b01111_011000_01111;
        tomato_rice_dim[29][5] = 16'b01111_011000_01111;
        tomato_rice_dim[29][6] = 16'b01111_011000_01111;
        tomato_rice_dim[29][7] = 16'b01111_011000_01111;
        tomato_rice_dim[29][8] = 16'b01111_011000_01111;
        tomato_rice_dim[29][9] = 16'b01111_011000_01111;
        tomato_rice_dim[29][10] = 16'b01111_011000_01111;
        tomato_rice_dim[29][11] = 16'b01111_011000_01111;
        tomato_rice_dim[29][12] = 16'b01111_011000_01111;
        tomato_rice_dim[29][13] = 16'b01111_011000_01111;
        tomato_rice_dim[29][14] = 16'b01111_011000_01111;
        tomato_rice_dim[29][15] = 16'b01111_011000_01111;
        tomato_rice_dim[29][16] = 16'b01111_011000_01111;
        tomato_rice_dim[29][17] = 16'b01111_011000_01111;
        tomato_rice_dim[29][18] = 16'b01111_011000_01111;
        tomato_rice_dim[29][19] = 16'b01111_011000_01111;
        tomato_rice_dim[29][20] = 16'b01111_011000_01111;
        tomato_rice_dim[29][21] = 16'b01111_011000_01111;
        tomato_rice_dim[29][22] = 16'b01111_011000_01111;
        tomato_rice_dim[29][23] = 16'b01111_011000_01111;
        tomato_rice_dim[29][24] = 16'b01111_011000_01111;
        tomato_rice_dim[29][25] = 16'b01111_011000_01111;
        tomato_rice_dim[29][26] = 16'b01111_011000_01111;
        tomato_rice_dim[29][27] = 16'b01111_011000_01111;
        tomato_rice_dim[29][28] = 16'b01111_011000_01111;
        tomato_rice_dim[29][29] = 16'b01111_011000_01111;
        tomato_rice_dim[29][30] = 16'b01111_011000_01111;
        tomato_rice_dim[29][31] = 16'b01111_011000_01111;
        tomato_rice_dim[30][0] = 16'b01111_011000_01111;
        tomato_rice_dim[30][1] = 16'b01111_011000_01111;
        tomato_rice_dim[30][2] = 16'b01111_011000_01111;
        tomato_rice_dim[30][3] = 16'b01111_011000_01111;
        tomato_rice_dim[30][4] = 16'b01111_011000_01111;
        tomato_rice_dim[30][5] = 16'b01111_011000_01111;
        tomato_rice_dim[30][6] = 16'b01111_011000_01111;
        tomato_rice_dim[30][7] = 16'b01111_011000_01111;
        tomato_rice_dim[30][8] = 16'b01111_011000_01111;
        tomato_rice_dim[30][9] = 16'b01111_011000_01111;
        tomato_rice_dim[30][10] = 16'b01111_011000_01111;
        tomato_rice_dim[30][11] = 16'b01111_011000_01111;
        tomato_rice_dim[30][12] = 16'b01111_011000_01111;
        tomato_rice_dim[30][13] = 16'b01111_011000_01111;
        tomato_rice_dim[30][14] = 16'b01111_011000_01111;
        tomato_rice_dim[30][15] = 16'b01111_011000_01111;
        tomato_rice_dim[30][16] = 16'b01111_011000_01111;
        tomato_rice_dim[30][17] = 16'b01111_011000_01111;
        tomato_rice_dim[30][18] = 16'b01111_011000_01111;
        tomato_rice_dim[30][19] = 16'b01111_011000_01111;
        tomato_rice_dim[30][20] = 16'b01111_011000_01111;
        tomato_rice_dim[30][21] = 16'b01111_011000_01111;
        tomato_rice_dim[30][22] = 16'b01111_011000_01111;
        tomato_rice_dim[30][23] = 16'b01111_011000_01111;
        tomato_rice_dim[30][24] = 16'b01111_011000_01111;
        tomato_rice_dim[30][25] = 16'b01111_011000_01111;
        tomato_rice_dim[30][26] = 16'b01111_011000_01111;
        tomato_rice_dim[30][27] = 16'b01111_011000_01111;
        tomato_rice_dim[30][28] = 16'b01111_011000_01111;
        tomato_rice_dim[30][29] = 16'b01111_011000_01111;
        tomato_rice_dim[30][30] = 16'b01111_011000_01111;
        tomato_rice_dim[30][31] = 16'b01111_011000_01111;
        tomato_rice_dim[31][0] = 16'b01111_011000_01111;
        tomato_rice_dim[31][1] = 16'b01111_011000_01111;
        tomato_rice_dim[31][2] = 16'b01111_011000_01111;
        tomato_rice_dim[31][3] = 16'b01111_011000_01111;
        tomato_rice_dim[31][4] = 16'b01111_011000_01111;
        tomato_rice_dim[31][5] = 16'b01111_011000_01111;
        tomato_rice_dim[31][6] = 16'b01111_011000_01111;
        tomato_rice_dim[31][7] = 16'b01111_011000_01111;
        tomato_rice_dim[31][8] = 16'b01111_011000_01111;
        tomato_rice_dim[31][9] = 16'b01111_011000_01111;
        tomato_rice_dim[31][10] = 16'b01111_011000_01111;
        tomato_rice_dim[31][11] = 16'b01111_011000_01111;
        tomato_rice_dim[31][12] = 16'b01111_011000_01111;
        tomato_rice_dim[31][13] = 16'b01111_011000_01111;
        tomato_rice_dim[31][14] = 16'b01111_011000_01111;
        tomato_rice_dim[31][15] = 16'b01111_011000_01111;
        tomato_rice_dim[31][16] = 16'b01111_011000_01111;
        tomato_rice_dim[31][17] = 16'b01111_011000_01111;
        tomato_rice_dim[31][18] = 16'b01111_011000_01111;
        tomato_rice_dim[31][19] = 16'b01111_011000_01111;
        tomato_rice_dim[31][20] = 16'b01111_011000_01111;
        tomato_rice_dim[31][21] = 16'b01111_011000_01111;
        tomato_rice_dim[31][22] = 16'b01111_011000_01111;
        tomato_rice_dim[31][23] = 16'b01111_011000_01111;
        tomato_rice_dim[31][24] = 16'b01111_011000_01111;
        tomato_rice_dim[31][25] = 16'b01111_011000_01111;
        tomato_rice_dim[31][26] = 16'b01111_011000_01111;
        tomato_rice_dim[31][27] = 16'b01111_011000_01111;
        tomato_rice_dim[31][28] = 16'b01111_011000_01111;
        tomato_rice_dim[31][29] = 16'b01111_011000_01111;
        tomato_rice_dim[31][30] = 16'b01111_011000_01111;
        tomato_rice_dim[31][31] = 16'b01111_011000_01111;


        
        ingredient_text[0][0] = 16'b00011_000110_00011;
        ingredient_text[0][1] = 16'b00011_000110_00011;
        ingredient_text[0][2] = 16'b00011_000110_00011;
        ingredient_text[0][3] = 16'b00011_000110_00011;
        ingredient_text[0][4] = 16'b00011_000110_00011;
        ingredient_text[0][5] = 16'b00011_000110_00011;
        ingredient_text[0][6] = 16'b00011_000110_00011;
        ingredient_text[0][7] = 16'b00011_000110_00011;
        ingredient_text[0][8] = 16'b00011_000110_00011;
        ingredient_text[0][9] = 16'b00011_000110_00011;
        ingredient_text[0][10] = 16'b00011_000110_00011;
        ingredient_text[0][11] = 16'b00011_000110_00011;
        ingredient_text[0][12] = 16'b00011_000110_00011;
        ingredient_text[0][13] = 16'b00011_000110_00011;
        ingredient_text[0][14] = 16'b00011_000110_00011;
        ingredient_text[0][15] = 16'b00011_000110_00011;
        ingredient_text[0][16] = 16'b00011_000110_00011;
        ingredient_text[0][17] = 16'b00011_000110_00011;
        ingredient_text[0][18] = 16'b00011_000110_00011;
        ingredient_text[0][19] = 16'b00011_000110_00011;
        ingredient_text[0][20] = 16'b00011_000110_00011;
        ingredient_text[0][21] = 16'b00011_000110_00011;
        ingredient_text[0][22] = 16'b00011_000110_00011;
        ingredient_text[0][23] = 16'b00011_000110_00011;
        ingredient_text[0][24] = 16'b00011_000110_00011;
        ingredient_text[0][25] = 16'b00011_000110_00011;
        ingredient_text[0][26] = 16'b00011_000110_00011;
        ingredient_text[0][27] = 16'b00011_000110_00011;
        ingredient_text[0][28] = 16'b00011_000110_00011;
        ingredient_text[0][29] = 16'b00011_000110_00011;
        ingredient_text[0][30] = 16'b00011_000110_00011;
        ingredient_text[0][31] = 16'b00011_000110_00011;
        ingredient_text[0][32] = 16'b00011_000110_00011;
        ingredient_text[0][33] = 16'b00011_000110_00011;
        ingredient_text[0][34] = 16'b00011_000110_00011;
        ingredient_text[0][35] = 16'b00011_000110_00011;
        ingredient_text[0][36] = 16'b00011_000110_00011;
        ingredient_text[0][37] = 16'b00011_000110_00011;
        ingredient_text[0][38] = 16'b00011_000110_00011;
        ingredient_text[0][39] = 16'b00011_000110_00011;
        ingredient_text[0][40] = 16'b00011_000110_00011;
        ingredient_text[0][41] = 16'b00011_000110_00011;
        ingredient_text[0][42] = 16'b00011_000110_00011;
        ingredient_text[0][43] = 16'b00011_000110_00011;
        ingredient_text[0][44] = 16'b00011_000110_00011;
        ingredient_text[0][45] = 16'b00011_000110_00011;
        ingredient_text[0][46] = 16'b00011_000110_00011;
        ingredient_text[0][47] = 16'b00011_000110_00011;
        ingredient_text[0][48] = 16'b00011_000110_00011;
        ingredient_text[0][49] = 16'b00011_000110_00011;
        ingredient_text[0][50] = 16'b00011_000110_00011;
        ingredient_text[0][51] = 16'b00011_000110_00011;
        ingredient_text[0][52] = 16'b00011_000110_00011;
        ingredient_text[0][53] = 16'b00011_000110_00011;
        ingredient_text[0][54] = 16'b00011_000110_00011;
        ingredient_text[0][55] = 16'b00011_000110_00011;
        ingredient_text[0][56] = 16'b00011_000110_00011;
        ingredient_text[0][57] = 16'b00011_000110_00011;
        ingredient_text[0][58] = 16'b00011_000110_00011;
        ingredient_text[0][59] = 16'b00011_000110_00011;
        ingredient_text[0][60] = 16'b00011_000110_00011;
        ingredient_text[0][61] = 16'b00011_000110_00011;
        ingredient_text[0][62] = 16'b00011_000110_00011;
        ingredient_text[0][63] = 16'b00011_000110_00011;
        ingredient_text[0][64] = 16'b00011_000110_00011;
        ingredient_text[0][65] = 16'b00011_000110_00011;
        ingredient_text[0][66] = 16'b00011_000110_00011;
        ingredient_text[0][67] = 16'b00011_000110_00011;
        ingredient_text[0][68] = 16'b00011_000110_00011;
        ingredient_text[0][69] = 16'b00011_000110_00011;
        ingredient_text[0][70] = 16'b00011_000110_00011;
        ingredient_text[0][71] = 16'b00011_000110_00011;
        ingredient_text[0][72] = 16'b00011_000110_00011;
        ingredient_text[0][73] = 16'b00011_000110_00011;
        ingredient_text[0][74] = 16'b00011_000110_00011;
        ingredient_text[0][75] = 16'b00011_000110_00011;
        ingredient_text[0][76] = 16'b00011_000110_00011;
        ingredient_text[0][77] = 16'b00011_000110_00011;
        ingredient_text[0][78] = 16'b00011_000110_00011;
        ingredient_text[0][79] = 16'b00011_000110_00011;
        ingredient_text[1][0] = 16'b00011_000110_00011;
        ingredient_text[1][1] = 16'b00011_000110_00011;
        ingredient_text[1][2] = 16'b00011_000110_00011;
        ingredient_text[1][3] = 16'b00011_000110_00011;
        ingredient_text[1][4] = 16'b00011_000110_00011;
        ingredient_text[1][5] = 16'b00011_000110_00011;
        ingredient_text[1][6] = 16'b00011_000110_00011;
        ingredient_text[1][7] = 16'b00011_000110_00011;
        ingredient_text[1][8] = 16'b00011_000110_00011;
        ingredient_text[1][9] = 16'b00011_000110_00011;
        ingredient_text[1][10] = 16'b00011_000110_00011;
        ingredient_text[1][11] = 16'b00011_000110_00011;
        ingredient_text[1][12] = 16'b00011_000110_00011;
        ingredient_text[1][13] = 16'b00011_000110_00011;
        ingredient_text[1][14] = 16'b00011_000110_00011;
        ingredient_text[1][15] = 16'b00011_000110_00011;
        ingredient_text[1][16] = 16'b00011_000110_00011;
        ingredient_text[1][17] = 16'b00011_000110_00011;
        ingredient_text[1][18] = 16'b00011_000110_00011;
        ingredient_text[1][19] = 16'b00011_000110_00011;
        ingredient_text[1][20] = 16'b00011_000110_00011;
        ingredient_text[1][21] = 16'b00011_000110_00011;
        ingredient_text[1][22] = 16'b00011_000110_00011;
        ingredient_text[1][23] = 16'b00011_000110_00011;
        ingredient_text[1][24] = 16'b00011_000110_00011;
        ingredient_text[1][25] = 16'b00011_000110_00011;
        ingredient_text[1][26] = 16'b00011_000110_00011;
        ingredient_text[1][27] = 16'b00011_000110_00011;
        ingredient_text[1][28] = 16'b00011_000110_00011;
        ingredient_text[1][29] = 16'b00011_000110_00011;
        ingredient_text[1][30] = 16'b00011_000110_00011;
        ingredient_text[1][31] = 16'b00011_000110_00011;
        ingredient_text[1][32] = 16'b00011_000110_00011;
        ingredient_text[1][33] = 16'b00011_000110_00011;
        ingredient_text[1][34] = 16'b00011_000110_00011;
        ingredient_text[1][35] = 16'b00011_000110_00011;
        ingredient_text[1][36] = 16'b00011_000110_00011;
        ingredient_text[1][37] = 16'b00011_000110_00011;
        ingredient_text[1][38] = 16'b00011_000110_00011;
        ingredient_text[1][39] = 16'b00011_000110_00011;
        ingredient_text[1][40] = 16'b00011_000110_00011;
        ingredient_text[1][41] = 16'b00011_000110_00011;
        ingredient_text[1][42] = 16'b00011_000110_00011;
        ingredient_text[1][43] = 16'b00011_000110_00011;
        ingredient_text[1][44] = 16'b00011_000110_00011;
        ingredient_text[1][45] = 16'b00011_000110_00011;
        ingredient_text[1][46] = 16'b00011_000110_00011;
        ingredient_text[1][47] = 16'b00011_000110_00011;
        ingredient_text[1][48] = 16'b00011_000110_00011;
        ingredient_text[1][49] = 16'b00011_000110_00011;
        ingredient_text[1][50] = 16'b00011_000110_00011;
        ingredient_text[1][51] = 16'b00011_000110_00011;
        ingredient_text[1][52] = 16'b00011_000110_00011;
        ingredient_text[1][53] = 16'b00011_000110_00011;
        ingredient_text[1][54] = 16'b00011_000110_00011;
        ingredient_text[1][55] = 16'b00011_000110_00011;
        ingredient_text[1][56] = 16'b00011_000110_00011;
        ingredient_text[1][57] = 16'b00011_000110_00011;
        ingredient_text[1][58] = 16'b00011_000110_00011;
        ingredient_text[1][59] = 16'b01110_011110_01110;
        ingredient_text[1][60] = 16'b11111_111111_11111;
        ingredient_text[1][61] = 16'b11111_111111_11111;
        ingredient_text[1][62] = 16'b11011_110111_11011;
        ingredient_text[1][63] = 16'b10110_101101_10110;
        ingredient_text[1][64] = 16'b00011_000110_00011;
        ingredient_text[1][65] = 16'b00011_000110_00011;
        ingredient_text[1][66] = 16'b00011_000110_00011;
        ingredient_text[1][67] = 16'b00011_000110_00011;
        ingredient_text[1][68] = 16'b00011_000110_00011;
        ingredient_text[1][69] = 16'b00011_000110_00011;
        ingredient_text[1][70] = 16'b00011_000110_00011;
        ingredient_text[1][71] = 16'b00011_000110_00011;
        ingredient_text[1][72] = 16'b00011_000110_00011;
        ingredient_text[1][73] = 16'b00011_000110_00011;
        ingredient_text[1][74] = 16'b00011_000110_00011;
        ingredient_text[1][75] = 16'b00011_000110_00011;
        ingredient_text[1][76] = 16'b00011_000110_00011;
        ingredient_text[1][77] = 16'b00011_000110_00011;
        ingredient_text[1][78] = 16'b00011_000110_00011;
        ingredient_text[1][79] = 16'b00011_000110_00011;
        ingredient_text[2][0] = 16'b00011_000110_00011;
        ingredient_text[2][1] = 16'b00011_000110_00011;
        ingredient_text[2][2] = 16'b00011_000110_00011;
        ingredient_text[2][3] = 16'b00011_000110_00011;
        ingredient_text[2][4] = 16'b00011_000110_00011;
        ingredient_text[2][5] = 16'b00011_000110_00011;
        ingredient_text[2][6] = 16'b00011_000110_00011;
        ingredient_text[2][7] = 16'b00011_000110_00011;
        ingredient_text[2][8] = 16'b00011_000110_00011;
        ingredient_text[2][9] = 16'b00011_000110_00011;
        ingredient_text[2][10] = 16'b00011_000110_00011;
        ingredient_text[2][11] = 16'b00011_000110_00011;
        ingredient_text[2][12] = 16'b00011_000110_00011;
        ingredient_text[2][13] = 16'b00011_000110_00011;
        ingredient_text[2][14] = 16'b00011_000110_00011;
        ingredient_text[2][15] = 16'b00011_000110_00011;
        ingredient_text[2][16] = 16'b00011_000110_00011;
        ingredient_text[2][17] = 16'b00011_000110_00011;
        ingredient_text[2][18] = 16'b00011_000110_00011;
        ingredient_text[2][19] = 16'b00011_000110_00011;
        ingredient_text[2][20] = 16'b00011_000110_00011;
        ingredient_text[2][21] = 16'b00011_000110_00011;
        ingredient_text[2][22] = 16'b00011_000110_00011;
        ingredient_text[2][23] = 16'b00011_000110_00011;
        ingredient_text[2][24] = 16'b00011_000110_00011;
        ingredient_text[2][25] = 16'b00011_000110_00011;
        ingredient_text[2][26] = 16'b00011_000110_00011;
        ingredient_text[2][27] = 16'b00011_000110_00011;
        ingredient_text[2][28] = 16'b00011_000110_00011;
        ingredient_text[2][29] = 16'b00011_000110_00011;
        ingredient_text[2][30] = 16'b00011_000110_00011;
        ingredient_text[2][31] = 16'b00011_000110_00011;
        ingredient_text[2][32] = 16'b00011_000110_00011;
        ingredient_text[2][33] = 16'b00011_000110_00011;
        ingredient_text[2][34] = 16'b00011_000110_00011;
        ingredient_text[2][35] = 16'b00011_000110_00011;
        ingredient_text[2][36] = 16'b00011_000110_00011;
        ingredient_text[2][37] = 16'b00011_000110_00011;
        ingredient_text[2][38] = 16'b00011_000110_00011;
        ingredient_text[2][39] = 16'b00011_000110_00011;
        ingredient_text[2][40] = 16'b00011_000110_00011;
        ingredient_text[2][41] = 16'b00011_000110_00011;
        ingredient_text[2][42] = 16'b00011_000110_00011;
        ingredient_text[2][43] = 16'b00011_000110_00011;
        ingredient_text[2][44] = 16'b00011_000110_00011;
        ingredient_text[2][45] = 16'b00011_000110_00011;
        ingredient_text[2][46] = 16'b00011_000110_00011;
        ingredient_text[2][47] = 16'b00011_000110_00011;
        ingredient_text[2][48] = 16'b00011_000110_00011;
        ingredient_text[2][49] = 16'b00011_000110_00011;
        ingredient_text[2][50] = 16'b00011_000110_00011;
        ingredient_text[2][51] = 16'b00011_000110_00011;
        ingredient_text[2][52] = 16'b00011_000110_00011;
        ingredient_text[2][53] = 16'b00011_000110_00011;
        ingredient_text[2][54] = 16'b00011_000110_00011;
        ingredient_text[2][55] = 16'b00011_000110_00011;
        ingredient_text[2][56] = 16'b00011_000110_00011;
        ingredient_text[2][57] = 16'b00011_000110_00011;
        ingredient_text[2][58] = 16'b01110_011110_01110;
        ingredient_text[2][59] = 16'b11111_111111_11111;
        ingredient_text[2][60] = 16'b11111_111111_11111;
        ingredient_text[2][61] = 16'b11111_111111_11111;
        ingredient_text[2][62] = 16'b11111_111111_11111;
        ingredient_text[2][63] = 16'b11111_111111_11111;
        ingredient_text[2][64] = 16'b01110_011110_01110;
        ingredient_text[2][65] = 16'b00011_000110_00011;
        ingredient_text[2][66] = 16'b00011_000110_00011;
        ingredient_text[2][67] = 16'b00011_000110_00011;
        ingredient_text[2][68] = 16'b00011_000110_00011;
        ingredient_text[2][69] = 16'b00011_000110_00011;
        ingredient_text[2][70] = 16'b00011_000110_00011;
        ingredient_text[2][71] = 16'b00011_000110_00011;
        ingredient_text[2][72] = 16'b00011_000110_00011;
        ingredient_text[2][73] = 16'b00011_000110_00011;
        ingredient_text[2][74] = 16'b00011_000110_00011;
        ingredient_text[2][75] = 16'b00011_000110_00011;
        ingredient_text[2][76] = 16'b00011_000110_00011;
        ingredient_text[2][77] = 16'b00011_000110_00011;
        ingredient_text[2][78] = 16'b00011_000110_00011;
        ingredient_text[2][79] = 16'b00011_000110_00011;
        ingredient_text[3][0] = 16'b00011_000110_00011;
        ingredient_text[3][1] = 16'b00011_000110_00011;
        ingredient_text[3][2] = 16'b00011_000110_00011;
        ingredient_text[3][3] = 16'b00011_000110_00011;
        ingredient_text[3][4] = 16'b00011_000110_00011;
        ingredient_text[3][5] = 16'b00011_000110_00011;
        ingredient_text[3][6] = 16'b00011_000110_00011;
        ingredient_text[3][7] = 16'b00011_000110_00011;
        ingredient_text[3][8] = 16'b00011_000110_00011;
        ingredient_text[3][9] = 16'b00011_000110_00011;
        ingredient_text[3][10] = 16'b00011_000110_00011;
        ingredient_text[3][11] = 16'b00011_000110_00011;
        ingredient_text[3][12] = 16'b00011_000110_00011;
        ingredient_text[3][13] = 16'b00011_000110_00011;
        ingredient_text[3][14] = 16'b00011_000110_00011;
        ingredient_text[3][15] = 16'b00011_000110_00011;
        ingredient_text[3][16] = 16'b00011_000110_00011;
        ingredient_text[3][17] = 16'b00011_000110_00011;
        ingredient_text[3][18] = 16'b00011_000110_00011;
        ingredient_text[3][19] = 16'b00011_000110_00011;
        ingredient_text[3][20] = 16'b00011_000110_00011;
        ingredient_text[3][21] = 16'b00011_000110_00011;
        ingredient_text[3][22] = 16'b00011_000110_00011;
        ingredient_text[3][23] = 16'b00011_000110_00011;
        ingredient_text[3][24] = 16'b00011_000110_00011;
        ingredient_text[3][25] = 16'b00011_000110_00011;
        ingredient_text[3][26] = 16'b00011_000110_00011;
        ingredient_text[3][27] = 16'b00011_000110_00011;
        ingredient_text[3][28] = 16'b00011_000110_00011;
        ingredient_text[3][29] = 16'b00011_000110_00011;
        ingredient_text[3][30] = 16'b00011_000110_00011;
        ingredient_text[3][31] = 16'b00011_000110_00011;
        ingredient_text[3][32] = 16'b00011_000110_00011;
        ingredient_text[3][33] = 16'b00011_000110_00011;
        ingredient_text[3][34] = 16'b00011_000110_00011;
        ingredient_text[3][35] = 16'b00011_000110_00011;
        ingredient_text[3][36] = 16'b00011_000110_00011;
        ingredient_text[3][37] = 16'b00011_000110_00011;
        ingredient_text[3][38] = 16'b00011_000110_00011;
        ingredient_text[3][39] = 16'b00011_000110_00011;
        ingredient_text[3][40] = 16'b00011_000110_00011;
        ingredient_text[3][41] = 16'b00011_000110_00011;
        ingredient_text[3][42] = 16'b00011_000110_00011;
        ingredient_text[3][43] = 16'b00011_000110_00011;
        ingredient_text[3][44] = 16'b00011_000110_00011;
        ingredient_text[3][45] = 16'b00011_000110_00011;
        ingredient_text[3][46] = 16'b00011_000110_00011;
        ingredient_text[3][47] = 16'b00011_000110_00011;
        ingredient_text[3][48] = 16'b00011_000110_00011;
        ingredient_text[3][49] = 16'b00011_000110_00011;
        ingredient_text[3][50] = 16'b00011_000110_00011;
        ingredient_text[3][51] = 16'b00011_000110_00011;
        ingredient_text[3][52] = 16'b00011_000110_00011;
        ingredient_text[3][53] = 16'b00011_000110_00011;
        ingredient_text[3][54] = 16'b00011_000110_00011;
        ingredient_text[3][55] = 16'b00011_000110_00011;
        ingredient_text[3][56] = 16'b00011_000110_00011;
        ingredient_text[3][57] = 16'b00011_000110_00011;
        ingredient_text[3][58] = 16'b11011_110111_11011;
        ingredient_text[3][59] = 16'b11111_111111_11111;
        ingredient_text[3][60] = 16'b00011_000110_00011;
        ingredient_text[3][61] = 16'b00011_000110_00011;
        ingredient_text[3][62] = 16'b01110_011110_01110;
        ingredient_text[3][63] = 16'b11111_111111_11111;
        ingredient_text[3][64] = 16'b01110_011110_01110;
        ingredient_text[3][65] = 16'b00011_000110_00011;
        ingredient_text[3][66] = 16'b00011_000110_00011;
        ingredient_text[3][67] = 16'b00011_000110_00011;
        ingredient_text[3][68] = 16'b00011_000110_00011;
        ingredient_text[3][69] = 16'b00011_000110_00011;
        ingredient_text[3][70] = 16'b00011_000110_00011;
        ingredient_text[3][71] = 16'b00011_000110_00011;
        ingredient_text[3][72] = 16'b00011_000110_00011;
        ingredient_text[3][73] = 16'b00011_000110_00011;
        ingredient_text[3][74] = 16'b00011_000110_00011;
        ingredient_text[3][75] = 16'b00011_000110_00011;
        ingredient_text[3][76] = 16'b00011_000110_00011;
        ingredient_text[3][77] = 16'b00011_000110_00011;
        ingredient_text[3][78] = 16'b00011_000110_00011;
        ingredient_text[3][79] = 16'b00011_000110_00011;
        ingredient_text[4][0] = 16'b00011_000110_00011;
        ingredient_text[4][1] = 16'b00011_000110_00011;
        ingredient_text[4][2] = 16'b00011_000110_00011;
        ingredient_text[4][3] = 16'b00011_000110_00011;
        ingredient_text[4][4] = 16'b00011_000110_00011;
        ingredient_text[4][5] = 16'b00011_000110_00011;
        ingredient_text[4][6] = 16'b00011_000110_00011;
        ingredient_text[4][7] = 16'b00011_000110_00011;
        ingredient_text[4][8] = 16'b00011_000110_00011;
        ingredient_text[4][9] = 16'b00011_000110_00011;
        ingredient_text[4][10] = 16'b00011_000110_00011;
        ingredient_text[4][11] = 16'b00011_000110_00011;
        ingredient_text[4][12] = 16'b00011_000110_00011;
        ingredient_text[4][13] = 16'b00011_000110_00011;
        ingredient_text[4][14] = 16'b00011_000110_00011;
        ingredient_text[4][15] = 16'b00011_000110_00011;
        ingredient_text[4][16] = 16'b11111_111111_11111;
        ingredient_text[4][17] = 16'b11111_111111_11111;
        ingredient_text[4][18] = 16'b11111_111111_11111;
        ingredient_text[4][19] = 16'b00011_000110_00011;
        ingredient_text[4][20] = 16'b00011_000110_00011;
        ingredient_text[4][21] = 16'b11011_110111_11011;
        ingredient_text[4][22] = 16'b11111_111111_11111;
        ingredient_text[4][23] = 16'b00011_000110_00011;
        ingredient_text[4][24] = 16'b00011_000110_00011;
        ingredient_text[4][25] = 16'b10110_101101_10110;
        ingredient_text[4][26] = 16'b11111_111111_11111;
        ingredient_text[4][27] = 16'b00011_000110_00011;
        ingredient_text[4][28] = 16'b00011_000110_00011;
        ingredient_text[4][29] = 16'b11111_111111_11111;
        ingredient_text[4][30] = 16'b11111_111111_11111;
        ingredient_text[4][31] = 16'b11111_111111_11111;
        ingredient_text[4][32] = 16'b11111_111111_11111;
        ingredient_text[4][33] = 16'b11011_110111_11011;
        ingredient_text[4][34] = 16'b00011_000110_00011;
        ingredient_text[4][35] = 16'b00011_000110_00011;
        ingredient_text[4][36] = 16'b11111_111111_11111;
        ingredient_text[4][37] = 16'b11011_110111_11011;
        ingredient_text[4][38] = 16'b00011_000110_00011;
        ingredient_text[4][39] = 16'b11011_110111_11011;
        ingredient_text[4][40] = 16'b11111_111111_11111;
        ingredient_text[4][41] = 16'b11111_111111_11111;
        ingredient_text[4][42] = 16'b11111_111111_11111;
        ingredient_text[4][43] = 16'b11111_111111_11111;
        ingredient_text[4][44] = 16'b11011_110111_11011;
        ingredient_text[4][45] = 16'b00011_000110_00011;
        ingredient_text[4][46] = 16'b00011_000110_00011;
        ingredient_text[4][47] = 16'b11111_111111_11111;
        ingredient_text[4][48] = 16'b11111_111111_11111;
        ingredient_text[4][49] = 16'b11111_111111_11111;
        ingredient_text[4][50] = 16'b11111_111111_11111;
        ingredient_text[4][51] = 16'b11011_110111_11011;
        ingredient_text[4][52] = 16'b00011_000110_00011;
        ingredient_text[4][53] = 16'b00011_000110_00011;
        ingredient_text[4][54] = 16'b00011_000110_00011;
        ingredient_text[4][55] = 16'b11111_111111_11111;
        ingredient_text[4][56] = 16'b11111_111111_11111;
        ingredient_text[4][57] = 16'b00011_000110_00011;
        ingredient_text[4][58] = 16'b00011_000110_00011;
        ingredient_text[4][59] = 16'b11111_111111_11111;
        ingredient_text[4][60] = 16'b11111_111111_11111;
        ingredient_text[4][61] = 16'b11111_111111_11111;
        ingredient_text[4][62] = 16'b11111_111111_11111;
        ingredient_text[4][63] = 16'b11111_111111_11111;
        ingredient_text[4][64] = 16'b00011_000110_00011;
        ingredient_text[4][65] = 16'b11011_110111_11011;
        ingredient_text[4][66] = 16'b11111_111111_11111;
        ingredient_text[4][67] = 16'b00011_000110_00011;
        ingredient_text[4][68] = 16'b00011_000110_00011;
        ingredient_text[4][69] = 16'b10110_101101_10110;
        ingredient_text[4][70] = 16'b11111_111111_11111;
        ingredient_text[4][71] = 16'b00011_000110_00011;
        ingredient_text[4][72] = 16'b00011_000110_00011;
        ingredient_text[4][73] = 16'b11111_111111_11111;
        ingredient_text[4][74] = 16'b11111_111111_11111;
        ingredient_text[4][75] = 16'b00011_000110_00011;
        ingredient_text[4][76] = 16'b00011_000110_00011;
        ingredient_text[4][77] = 16'b00011_000110_00011;
        ingredient_text[4][78] = 16'b00011_000110_00011;
        ingredient_text[4][79] = 16'b00011_000110_00011;
        ingredient_text[5][0] = 16'b00011_000110_00011;
        ingredient_text[5][1] = 16'b00011_000110_00011;
        ingredient_text[5][2] = 16'b00011_000110_00011;
        ingredient_text[5][3] = 16'b00011_000110_00011;
        ingredient_text[5][4] = 16'b00011_000110_00011;
        ingredient_text[5][5] = 16'b00011_000110_00011;
        ingredient_text[5][6] = 16'b00011_000110_00011;
        ingredient_text[5][7] = 16'b00011_000110_00011;
        ingredient_text[5][8] = 16'b00011_000110_00011;
        ingredient_text[5][9] = 16'b00011_000110_00011;
        ingredient_text[5][10] = 16'b00011_000110_00011;
        ingredient_text[5][11] = 16'b00011_000110_00011;
        ingredient_text[5][12] = 16'b00011_000110_00011;
        ingredient_text[5][13] = 16'b00011_000110_00011;
        ingredient_text[5][14] = 16'b00011_000110_00011;
        ingredient_text[5][15] = 16'b00011_000110_00011;
        ingredient_text[5][16] = 16'b01110_011110_01110;
        ingredient_text[5][17] = 16'b01110_011110_01110;
        ingredient_text[5][18] = 16'b11111_111111_11111;
        ingredient_text[5][19] = 16'b10110_101101_10110;
        ingredient_text[5][20] = 16'b00011_000110_00011;
        ingredient_text[5][21] = 16'b11011_110111_11011;
        ingredient_text[5][22] = 16'b11111_111111_11111;
        ingredient_text[5][23] = 16'b00011_000110_00011;
        ingredient_text[5][24] = 16'b00011_000110_00011;
        ingredient_text[5][25] = 16'b10110_101101_10110;
        ingredient_text[5][26] = 16'b11111_111111_11111;
        ingredient_text[5][27] = 16'b00011_000110_00011;
        ingredient_text[5][28] = 16'b00011_000110_00011;
        ingredient_text[5][29] = 16'b10110_101101_10110;
        ingredient_text[5][30] = 16'b00011_000110_00011;
        ingredient_text[5][31] = 16'b00011_000110_00011;
        ingredient_text[5][32] = 16'b11011_110111_11011;
        ingredient_text[5][33] = 16'b11111_111111_11111;
        ingredient_text[5][34] = 16'b00011_000110_00011;
        ingredient_text[5][35] = 16'b00011_000110_00011;
        ingredient_text[5][36] = 16'b11111_111111_11111;
        ingredient_text[5][37] = 16'b11011_110111_11011;
        ingredient_text[5][38] = 16'b00011_000110_00011;
        ingredient_text[5][39] = 16'b11011_110111_11011;
        ingredient_text[5][40] = 16'b11111_111111_11111;
        ingredient_text[5][41] = 16'b11011_110111_11011;
        ingredient_text[5][42] = 16'b00011_000110_00011;
        ingredient_text[5][43] = 16'b11111_111111_11111;
        ingredient_text[5][44] = 16'b11111_111111_11111;
        ingredient_text[5][45] = 16'b00011_000110_00011;
        ingredient_text[5][46] = 16'b00011_000110_00011;
        ingredient_text[5][47] = 16'b10110_101101_10110;
        ingredient_text[5][48] = 16'b00011_000110_00011;
        ingredient_text[5][49] = 16'b00011_000110_00011;
        ingredient_text[5][50] = 16'b11011_110111_11011;
        ingredient_text[5][51] = 16'b11111_111111_11111;
        ingredient_text[5][52] = 16'b00011_000110_00011;
        ingredient_text[5][53] = 16'b00011_000110_00011;
        ingredient_text[5][54] = 16'b00011_000110_00011;
        ingredient_text[5][55] = 16'b11111_111111_11111;
        ingredient_text[5][56] = 16'b11111_111111_11111;
        ingredient_text[5][57] = 16'b00011_000110_00011;
        ingredient_text[5][58] = 16'b00011_000110_00011;
        ingredient_text[5][59] = 16'b00011_000110_00011;
        ingredient_text[5][60] = 16'b00011_000110_00011;
        ingredient_text[5][61] = 16'b00011_000110_00011;
        ingredient_text[5][62] = 16'b10110_101101_10110;
        ingredient_text[5][63] = 16'b11111_111111_11111;
        ingredient_text[5][64] = 16'b00011_000110_00011;
        ingredient_text[5][65] = 16'b11011_110111_11011;
        ingredient_text[5][66] = 16'b11111_111111_11111;
        ingredient_text[5][67] = 16'b00011_000110_00011;
        ingredient_text[5][68] = 16'b00011_000110_00011;
        ingredient_text[5][69] = 16'b10110_101101_10110;
        ingredient_text[5][70] = 16'b11111_111111_11111;
        ingredient_text[5][71] = 16'b00011_000110_00011;
        ingredient_text[5][72] = 16'b00011_000110_00011;
        ingredient_text[5][73] = 16'b11111_111111_11111;
        ingredient_text[5][74] = 16'b11111_111111_11111;
        ingredient_text[5][75] = 16'b00011_000110_00011;
        ingredient_text[5][76] = 16'b00011_000110_00011;
        ingredient_text[5][77] = 16'b00011_000110_00011;
        ingredient_text[5][78] = 16'b00011_000110_00011;
        ingredient_text[5][79] = 16'b00011_000110_00011;
        ingredient_text[6][0] = 16'b00011_000110_00011;
        ingredient_text[6][1] = 16'b00011_000110_00011;
        ingredient_text[6][2] = 16'b00011_000110_00011;
        ingredient_text[6][3] = 16'b00011_000110_00011;
        ingredient_text[6][4] = 16'b00011_000110_00011;
        ingredient_text[6][5] = 16'b00011_000110_00011;
        ingredient_text[6][6] = 16'b00011_000110_00011;
        ingredient_text[6][7] = 16'b00011_000110_00011;
        ingredient_text[6][8] = 16'b00011_000110_00011;
        ingredient_text[6][9] = 16'b00011_000110_00011;
        ingredient_text[6][10] = 16'b00011_000110_00011;
        ingredient_text[6][11] = 16'b00011_000110_00011;
        ingredient_text[6][12] = 16'b00011_000110_00011;
        ingredient_text[6][13] = 16'b00011_000110_00011;
        ingredient_text[6][14] = 16'b00011_000110_00011;
        ingredient_text[6][15] = 16'b00011_000110_00011;
        ingredient_text[6][16] = 16'b00011_000110_00011;
        ingredient_text[6][17] = 16'b00011_000110_00011;
        ingredient_text[6][18] = 16'b11111_111111_11111;
        ingredient_text[6][19] = 16'b10110_101101_10110;
        ingredient_text[6][20] = 16'b00011_000110_00011;
        ingredient_text[6][21] = 16'b11011_110111_11011;
        ingredient_text[6][22] = 16'b11111_111111_11111;
        ingredient_text[6][23] = 16'b00011_000110_00011;
        ingredient_text[6][24] = 16'b00011_000110_00011;
        ingredient_text[6][25] = 16'b10110_101101_10110;
        ingredient_text[6][26] = 16'b11111_111111_11111;
        ingredient_text[6][27] = 16'b00011_000110_00011;
        ingredient_text[6][28] = 16'b01110_011110_01110;
        ingredient_text[6][29] = 16'b11111_111111_11111;
        ingredient_text[6][30] = 16'b11111_111111_11111;
        ingredient_text[6][31] = 16'b11111_111111_11111;
        ingredient_text[6][32] = 16'b11111_111111_11111;
        ingredient_text[6][33] = 16'b11111_111111_11111;
        ingredient_text[6][34] = 16'b10110_101101_10110;
        ingredient_text[6][35] = 16'b00011_000110_00011;
        ingredient_text[6][36] = 16'b11111_111111_11111;
        ingredient_text[6][37] = 16'b11011_110111_11011;
        ingredient_text[6][38] = 16'b00011_000110_00011;
        ingredient_text[6][39] = 16'b11011_110111_11011;
        ingredient_text[6][40] = 16'b11111_111111_11111;
        ingredient_text[6][41] = 16'b00011_000110_00011;
        ingredient_text[6][42] = 16'b00011_000110_00011;
        ingredient_text[6][43] = 16'b00011_000110_00011;
        ingredient_text[6][44] = 16'b11111_111111_11111;
        ingredient_text[6][45] = 16'b10110_101101_10110;
        ingredient_text[6][46] = 16'b01110_011110_01110;
        ingredient_text[6][47] = 16'b11111_111111_11111;
        ingredient_text[6][48] = 16'b11111_111111_11111;
        ingredient_text[6][49] = 16'b11111_111111_11111;
        ingredient_text[6][50] = 16'b11111_111111_11111;
        ingredient_text[6][51] = 16'b11111_111111_11111;
        ingredient_text[6][52] = 16'b10110_101101_10110;
        ingredient_text[6][53] = 16'b00011_000110_00011;
        ingredient_text[6][54] = 16'b00011_000110_00011;
        ingredient_text[6][55] = 16'b11111_111111_11111;
        ingredient_text[6][56] = 16'b11111_111111_11111;
        ingredient_text[6][57] = 16'b00011_000110_00011;
        ingredient_text[6][58] = 16'b00011_000110_00011;
        ingredient_text[6][59] = 16'b10110_101101_10110;
        ingredient_text[6][60] = 16'b11111_111111_11111;
        ingredient_text[6][61] = 16'b11111_111111_11111;
        ingredient_text[6][62] = 16'b11111_111111_11111;
        ingredient_text[6][63] = 16'b11011_110111_11011;
        ingredient_text[6][64] = 16'b00011_000110_00011;
        ingredient_text[6][65] = 16'b11011_110111_11011;
        ingredient_text[6][66] = 16'b11111_111111_11111;
        ingredient_text[6][67] = 16'b00011_000110_00011;
        ingredient_text[6][68] = 16'b00011_000110_00011;
        ingredient_text[6][69] = 16'b10110_101101_10110;
        ingredient_text[6][70] = 16'b11111_111111_11111;
        ingredient_text[6][71] = 16'b00011_000110_00011;
        ingredient_text[6][72] = 16'b00011_000110_00011;
        ingredient_text[6][73] = 16'b11111_111111_11111;
        ingredient_text[6][74] = 16'b11111_111111_11111;
        ingredient_text[6][75] = 16'b00011_000110_00011;
        ingredient_text[6][76] = 16'b00011_000110_00011;
        ingredient_text[6][77] = 16'b00011_000110_00011;
        ingredient_text[6][78] = 16'b00011_000110_00011;
        ingredient_text[6][79] = 16'b00011_000110_00011;
        ingredient_text[7][0] = 16'b00011_000110_00011;
        ingredient_text[7][1] = 16'b00011_000110_00011;
        ingredient_text[7][2] = 16'b00011_000110_00011;
        ingredient_text[7][3] = 16'b00011_000110_00011;
        ingredient_text[7][4] = 16'b00011_000110_00011;
        ingredient_text[7][5] = 16'b00011_000110_00011;
        ingredient_text[7][6] = 16'b00011_000110_00011;
        ingredient_text[7][7] = 16'b00011_000110_00011;
        ingredient_text[7][8] = 16'b00011_000110_00011;
        ingredient_text[7][9] = 16'b00011_000110_00011;
        ingredient_text[7][10] = 16'b00011_000110_00011;
        ingredient_text[7][11] = 16'b00011_000110_00011;
        ingredient_text[7][12] = 16'b00011_000110_00011;
        ingredient_text[7][13] = 16'b00011_000110_00011;
        ingredient_text[7][14] = 16'b00011_000110_00011;
        ingredient_text[7][15] = 16'b00011_000110_00011;
        ingredient_text[7][16] = 16'b00011_000110_00011;
        ingredient_text[7][17] = 16'b00011_000110_00011;
        ingredient_text[7][18] = 16'b11111_111111_11111;
        ingredient_text[7][19] = 16'b10110_101101_10110;
        ingredient_text[7][20] = 16'b00011_000110_00011;
        ingredient_text[7][21] = 16'b11011_110111_11011;
        ingredient_text[7][22] = 16'b11111_111111_11111;
        ingredient_text[7][23] = 16'b00011_000110_00011;
        ingredient_text[7][24] = 16'b00011_000110_00011;
        ingredient_text[7][25] = 16'b10110_101101_10110;
        ingredient_text[7][26] = 16'b11111_111111_11111;
        ingredient_text[7][27] = 16'b00011_000110_00011;
        ingredient_text[7][28] = 16'b10110_101101_10110;
        ingredient_text[7][29] = 16'b11111_111111_11111;
        ingredient_text[7][30] = 16'b10110_101101_10110;
        ingredient_text[7][31] = 16'b10110_101101_10110;
        ingredient_text[7][32] = 16'b10110_101101_10110;
        ingredient_text[7][33] = 16'b11111_111111_11111;
        ingredient_text[7][34] = 16'b10110_101101_10110;
        ingredient_text[7][35] = 16'b00011_000110_00011;
        ingredient_text[7][36] = 16'b11111_111111_11111;
        ingredient_text[7][37] = 16'b11011_110111_11011;
        ingredient_text[7][38] = 16'b00011_000110_00011;
        ingredient_text[7][39] = 16'b11011_110111_11011;
        ingredient_text[7][40] = 16'b11111_111111_11111;
        ingredient_text[7][41] = 16'b00011_000110_00011;
        ingredient_text[7][42] = 16'b00011_000110_00011;
        ingredient_text[7][43] = 16'b01110_011110_01110;
        ingredient_text[7][44] = 16'b11111_111111_11111;
        ingredient_text[7][45] = 16'b01110_011110_01110;
        ingredient_text[7][46] = 16'b10110_101101_10110;
        ingredient_text[7][47] = 16'b11111_111111_11111;
        ingredient_text[7][48] = 16'b10110_101101_10110;
        ingredient_text[7][49] = 16'b10110_101101_10110;
        ingredient_text[7][50] = 16'b10110_101101_10110;
        ingredient_text[7][51] = 16'b11111_111111_11111;
        ingredient_text[7][52] = 16'b10110_101101_10110;
        ingredient_text[7][53] = 16'b00011_000110_00011;
        ingredient_text[7][54] = 16'b00011_000110_00011;
        ingredient_text[7][55] = 16'b11111_111111_11111;
        ingredient_text[7][56] = 16'b11111_111111_11111;
        ingredient_text[7][57] = 16'b00011_000110_00011;
        ingredient_text[7][58] = 16'b00011_000110_00011;
        ingredient_text[7][59] = 16'b11111_111111_11111;
        ingredient_text[7][60] = 16'b11011_110111_11011;
        ingredient_text[7][61] = 16'b00011_000110_00011;
        ingredient_text[7][62] = 16'b11011_110111_11011;
        ingredient_text[7][63] = 16'b11111_111111_11111;
        ingredient_text[7][64] = 16'b00011_000110_00011;
        ingredient_text[7][65] = 16'b11011_110111_11011;
        ingredient_text[7][66] = 16'b11111_111111_11111;
        ingredient_text[7][67] = 16'b00011_000110_00011;
        ingredient_text[7][68] = 16'b00011_000110_00011;
        ingredient_text[7][69] = 16'b10110_101101_10110;
        ingredient_text[7][70] = 16'b11111_111111_11111;
        ingredient_text[7][71] = 16'b00011_000110_00011;
        ingredient_text[7][72] = 16'b00011_000110_00011;
        ingredient_text[7][73] = 16'b11111_111111_11111;
        ingredient_text[7][74] = 16'b11111_111111_11111;
        ingredient_text[7][75] = 16'b00011_000110_00011;
        ingredient_text[7][76] = 16'b00011_000110_00011;
        ingredient_text[7][77] = 16'b00011_000110_00011;
        ingredient_text[7][78] = 16'b00011_000110_00011;
        ingredient_text[7][79] = 16'b00011_000110_00011;
        ingredient_text[8][0] = 16'b00011_000110_00011;
        ingredient_text[8][1] = 16'b00011_000110_00011;
        ingredient_text[8][2] = 16'b00011_000110_00011;
        ingredient_text[8][3] = 16'b00011_000110_00011;
        ingredient_text[8][4] = 16'b00011_000110_00011;
        ingredient_text[8][5] = 16'b00011_000110_00011;
        ingredient_text[8][6] = 16'b00011_000110_00011;
        ingredient_text[8][7] = 16'b00011_000110_00011;
        ingredient_text[8][8] = 16'b00011_000110_00011;
        ingredient_text[8][9] = 16'b00011_000110_00011;
        ingredient_text[8][10] = 16'b00011_000110_00011;
        ingredient_text[8][11] = 16'b00011_000110_00011;
        ingredient_text[8][12] = 16'b00011_000110_00011;
        ingredient_text[8][13] = 16'b00011_000110_00011;
        ingredient_text[8][14] = 16'b00011_000110_00011;
        ingredient_text[8][15] = 16'b00011_000110_00011;
        ingredient_text[8][16] = 16'b00011_000110_00011;
        ingredient_text[8][17] = 16'b00011_000110_00011;
        ingredient_text[8][18] = 16'b11111_111111_11111;
        ingredient_text[8][19] = 16'b10110_101101_10110;
        ingredient_text[8][20] = 16'b00011_000110_00011;
        ingredient_text[8][21] = 16'b10110_101101_10110;
        ingredient_text[8][22] = 16'b11111_111111_11111;
        ingredient_text[8][23] = 16'b11011_110111_11011;
        ingredient_text[8][24] = 16'b01110_011110_01110;
        ingredient_text[8][25] = 16'b11111_111111_11111;
        ingredient_text[8][26] = 16'b11111_111111_11111;
        ingredient_text[8][27] = 16'b00011_000110_00011;
        ingredient_text[8][28] = 16'b00011_000110_00011;
        ingredient_text[8][29] = 16'b11111_111111_11111;
        ingredient_text[8][30] = 16'b11011_110111_11011;
        ingredient_text[8][31] = 16'b00011_000110_00011;
        ingredient_text[8][32] = 16'b11011_110111_11011;
        ingredient_text[8][33] = 16'b11111_111111_11111;
        ingredient_text[8][34] = 16'b00011_000110_00011;
        ingredient_text[8][35] = 16'b00011_000110_00011;
        ingredient_text[8][36] = 16'b11111_111111_11111;
        ingredient_text[8][37] = 16'b11011_110111_11011;
        ingredient_text[8][38] = 16'b00011_000110_00011;
        ingredient_text[8][39] = 16'b11011_110111_11011;
        ingredient_text[8][40] = 16'b11111_111111_11111;
        ingredient_text[8][41] = 16'b11011_110111_11011;
        ingredient_text[8][42] = 16'b00011_000110_00011;
        ingredient_text[8][43] = 16'b11111_111111_11111;
        ingredient_text[8][44] = 16'b11111_111111_11111;
        ingredient_text[8][45] = 16'b00011_000110_00011;
        ingredient_text[8][46] = 16'b00011_000110_00011;
        ingredient_text[8][47] = 16'b11111_111111_11111;
        ingredient_text[8][48] = 16'b11011_110111_11011;
        ingredient_text[8][49] = 16'b00011_000110_00011;
        ingredient_text[8][50] = 16'b11011_110111_11011;
        ingredient_text[8][51] = 16'b11111_111111_11111;
        ingredient_text[8][52] = 16'b00011_000110_00011;
        ingredient_text[8][53] = 16'b01110_011110_01110;
        ingredient_text[8][54] = 16'b01110_011110_01110;
        ingredient_text[8][55] = 16'b11111_111111_11111;
        ingredient_text[8][56] = 16'b11111_111111_11111;
        ingredient_text[8][57] = 16'b00011_000110_00011;
        ingredient_text[8][58] = 16'b00011_000110_00011;
        ingredient_text[8][59] = 16'b11111_111111_11111;
        ingredient_text[8][60] = 16'b11011_110111_11011;
        ingredient_text[8][61] = 16'b00011_000110_00011;
        ingredient_text[8][62] = 16'b11011_110111_11011;
        ingredient_text[8][63] = 16'b11111_111111_11111;
        ingredient_text[8][64] = 16'b00011_000110_00011;
        ingredient_text[8][65] = 16'b10110_101101_10110;
        ingredient_text[8][66] = 16'b11111_111111_11111;
        ingredient_text[8][67] = 16'b11011_110111_11011;
        ingredient_text[8][68] = 16'b01110_011110_01110;
        ingredient_text[8][69] = 16'b11111_111111_11111;
        ingredient_text[8][70] = 16'b11111_111111_11111;
        ingredient_text[8][71] = 16'b00011_000110_00011;
        ingredient_text[8][72] = 16'b00011_000110_00011;
        ingredient_text[8][73] = 16'b11111_111111_11111;
        ingredient_text[8][74] = 16'b11111_111111_11111;
        ingredient_text[8][75] = 16'b00011_000110_00011;
        ingredient_text[8][76] = 16'b00011_000110_00011;
        ingredient_text[8][77] = 16'b00011_000110_00011;
        ingredient_text[8][78] = 16'b00011_000110_00011;
        ingredient_text[8][79] = 16'b00011_000110_00011;
        ingredient_text[9][0] = 16'b00011_000110_00011;
        ingredient_text[9][1] = 16'b00011_000110_00011;
        ingredient_text[9][2] = 16'b00011_000110_00011;
        ingredient_text[9][3] = 16'b00011_000110_00011;
        ingredient_text[9][4] = 16'b00011_000110_00011;
        ingredient_text[9][5] = 16'b00011_000110_00011;
        ingredient_text[9][6] = 16'b00011_000110_00011;
        ingredient_text[9][7] = 16'b00011_000110_00011;
        ingredient_text[9][8] = 16'b00011_000110_00011;
        ingredient_text[9][9] = 16'b00011_000110_00011;
        ingredient_text[9][10] = 16'b00011_000110_00011;
        ingredient_text[9][11] = 16'b00011_000110_00011;
        ingredient_text[9][12] = 16'b00011_000110_00011;
        ingredient_text[9][13] = 16'b00011_000110_00011;
        ingredient_text[9][14] = 16'b00011_000110_00011;
        ingredient_text[9][15] = 16'b00011_000110_00011;
        ingredient_text[9][16] = 16'b11111_111111_11111;
        ingredient_text[9][17] = 16'b11111_111111_11111;
        ingredient_text[9][18] = 16'b11111_111111_11111;
        ingredient_text[9][19] = 16'b11111_111111_11111;
        ingredient_text[9][20] = 16'b10110_101101_10110;
        ingredient_text[9][21] = 16'b00011_000110_00011;
        ingredient_text[9][22] = 16'b11111_111111_11111;
        ingredient_text[9][23] = 16'b11111_111111_11111;
        ingredient_text[9][24] = 16'b11111_111111_11111;
        ingredient_text[9][25] = 16'b10110_101101_10110;
        ingredient_text[9][26] = 16'b11111_111111_11111;
        ingredient_text[9][27] = 16'b00011_000110_00011;
        ingredient_text[9][28] = 16'b00011_000110_00011;
        ingredient_text[9][29] = 16'b11011_110111_11011;
        ingredient_text[9][30] = 16'b11111_111111_11111;
        ingredient_text[9][31] = 16'b11111_111111_11111;
        ingredient_text[9][32] = 16'b11111_111111_11111;
        ingredient_text[9][33] = 16'b10110_101101_10110;
        ingredient_text[9][34] = 16'b00011_000110_00011;
        ingredient_text[9][35] = 16'b00011_000110_00011;
        ingredient_text[9][36] = 16'b11111_111111_11111;
        ingredient_text[9][37] = 16'b11011_110111_11011;
        ingredient_text[9][38] = 16'b00011_000110_00011;
        ingredient_text[9][39] = 16'b11011_110111_11011;
        ingredient_text[9][40] = 16'b11111_111111_11111;
        ingredient_text[9][41] = 16'b11111_111111_11111;
        ingredient_text[9][42] = 16'b11111_111111_11111;
        ingredient_text[9][43] = 16'b11111_111111_11111;
        ingredient_text[9][44] = 16'b11011_110111_11011;
        ingredient_text[9][45] = 16'b00011_000110_00011;
        ingredient_text[9][46] = 16'b00011_000110_00011;
        ingredient_text[9][47] = 16'b11011_110111_11011;
        ingredient_text[9][48] = 16'b11111_111111_11111;
        ingredient_text[9][49] = 16'b11111_111111_11111;
        ingredient_text[9][50] = 16'b11111_111111_11111;
        ingredient_text[9][51] = 16'b10110_101101_10110;
        ingredient_text[9][52] = 16'b00011_000110_00011;
        ingredient_text[9][53] = 16'b11111_111111_11111;
        ingredient_text[9][54] = 16'b11111_111111_11111;
        ingredient_text[9][55] = 16'b11011_110111_11011;
        ingredient_text[9][56] = 16'b11111_111111_11111;
        ingredient_text[9][57] = 16'b00011_000110_00011;
        ingredient_text[9][58] = 16'b11111_111111_11111;
        ingredient_text[9][59] = 16'b11111_111111_11111;
        ingredient_text[9][60] = 16'b11111_111111_11111;
        ingredient_text[9][61] = 16'b11111_111111_11111;
        ingredient_text[9][62] = 16'b11111_111111_11111;
        ingredient_text[9][63] = 16'b01110_011110_01110;
        ingredient_text[9][64] = 16'b00011_000110_00011;
        ingredient_text[9][65] = 16'b00011_000110_00011;
        ingredient_text[9][66] = 16'b11111_111111_11111;
        ingredient_text[9][67] = 16'b11111_111111_11111;
        ingredient_text[9][68] = 16'b11111_111111_11111;
        ingredient_text[9][69] = 16'b10110_101101_10110;
        ingredient_text[9][70] = 16'b11111_111111_11111;
        ingredient_text[9][71] = 16'b00011_000110_00011;
        ingredient_text[9][72] = 16'b00011_000110_00011;
        ingredient_text[9][73] = 16'b11111_111111_11111;
        ingredient_text[9][74] = 16'b11111_111111_11111;
        ingredient_text[9][75] = 16'b00011_000110_00011;
        ingredient_text[9][76] = 16'b00011_000110_00011;
        ingredient_text[9][77] = 16'b00011_000110_00011;
        ingredient_text[9][78] = 16'b00011_000110_00011;
        ingredient_text[9][79] = 16'b00011_000110_00011;
        ingredient_text[10][0] = 16'b00011_000110_00011;
        ingredient_text[10][1] = 16'b00011_000110_00011;
        ingredient_text[10][2] = 16'b00011_000110_00011;
        ingredient_text[10][3] = 16'b00011_000110_00011;
        ingredient_text[10][4] = 16'b00011_000110_00011;
        ingredient_text[10][5] = 16'b00011_000110_00011;
        ingredient_text[10][6] = 16'b00011_000110_00011;
        ingredient_text[10][7] = 16'b00011_000110_00011;
        ingredient_text[10][8] = 16'b00011_000110_00011;
        ingredient_text[10][9] = 16'b00011_000110_00011;
        ingredient_text[10][10] = 16'b00011_000110_00011;
        ingredient_text[10][11] = 16'b00011_000110_00011;
        ingredient_text[10][12] = 16'b00011_000110_00011;
        ingredient_text[10][13] = 16'b00011_000110_00011;
        ingredient_text[10][14] = 16'b00011_000110_00011;
        ingredient_text[10][15] = 16'b00011_000110_00011;
        ingredient_text[10][16] = 16'b00011_000110_00011;
        ingredient_text[10][17] = 16'b00011_000110_00011;
        ingredient_text[10][18] = 16'b11111_111111_11111;
        ingredient_text[10][19] = 16'b10110_101101_10110;
        ingredient_text[10][20] = 16'b00011_000110_00011;
        ingredient_text[10][21] = 16'b00011_000110_00011;
        ingredient_text[10][22] = 16'b00011_000110_00011;
        ingredient_text[10][23] = 16'b00011_000110_00011;
        ingredient_text[10][24] = 16'b00011_000110_00011;
        ingredient_text[10][25] = 16'b00011_000110_00011;
        ingredient_text[10][26] = 16'b00011_000110_00011;
        ingredient_text[10][27] = 16'b00011_000110_00011;
        ingredient_text[10][28] = 16'b00011_000110_00011;
        ingredient_text[10][29] = 16'b00011_000110_00011;
        ingredient_text[10][30] = 16'b00011_000110_00011;
        ingredient_text[10][31] = 16'b00011_000110_00011;
        ingredient_text[10][32] = 16'b00011_000110_00011;
        ingredient_text[10][33] = 16'b00011_000110_00011;
        ingredient_text[10][34] = 16'b00011_000110_00011;
        ingredient_text[10][35] = 16'b00011_000110_00011;
        ingredient_text[10][36] = 16'b00011_000110_00011;
        ingredient_text[10][37] = 16'b00011_000110_00011;
        ingredient_text[10][38] = 16'b00011_000110_00011;
        ingredient_text[10][39] = 16'b11011_110111_11011;
        ingredient_text[10][40] = 16'b11111_111111_11111;
        ingredient_text[10][41] = 16'b00011_000110_00011;
        ingredient_text[10][42] = 16'b00011_000110_00011;
        ingredient_text[10][43] = 16'b00011_000110_00011;
        ingredient_text[10][44] = 16'b00011_000110_00011;
        ingredient_text[10][45] = 16'b00011_000110_00011;
        ingredient_text[10][46] = 16'b00011_000110_00011;
        ingredient_text[10][47] = 16'b00011_000110_00011;
        ingredient_text[10][48] = 16'b00011_000110_00011;
        ingredient_text[10][49] = 16'b00011_000110_00011;
        ingredient_text[10][50] = 16'b00011_000110_00011;
        ingredient_text[10][51] = 16'b00011_000110_00011;
        ingredient_text[10][52] = 16'b00011_000110_00011;
        ingredient_text[10][53] = 16'b00011_000110_00011;
        ingredient_text[10][54] = 16'b00011_000110_00011;
        ingredient_text[10][55] = 16'b00011_000110_00011;
        ingredient_text[10][56] = 16'b00011_000110_00011;
        ingredient_text[10][57] = 16'b00011_000110_00011;
        ingredient_text[10][58] = 16'b00011_000110_00011;
        ingredient_text[10][59] = 16'b00011_000110_00011;
        ingredient_text[10][60] = 16'b00011_000110_00011;
        ingredient_text[10][61] = 16'b00011_000110_00011;
        ingredient_text[10][62] = 16'b00011_000110_00011;
        ingredient_text[10][63] = 16'b00011_000110_00011;
        ingredient_text[10][64] = 16'b00011_000110_00011;
        ingredient_text[10][65] = 16'b00011_000110_00011;
        ingredient_text[10][66] = 16'b00011_000110_00011;
        ingredient_text[10][67] = 16'b00011_000110_00011;
        ingredient_text[10][68] = 16'b00011_000110_00011;
        ingredient_text[10][69] = 16'b00011_000110_00011;
        ingredient_text[10][70] = 16'b00011_000110_00011;
        ingredient_text[10][71] = 16'b00011_000110_00011;
        ingredient_text[10][72] = 16'b00011_000110_00011;
        ingredient_text[10][73] = 16'b11111_111111_11111;
        ingredient_text[10][74] = 16'b11111_111111_11111;
        ingredient_text[10][75] = 16'b00011_000110_00011;
        ingredient_text[10][76] = 16'b00011_000110_00011;
        ingredient_text[10][77] = 16'b00011_000110_00011;
        ingredient_text[10][78] = 16'b00011_000110_00011;
        ingredient_text[10][79] = 16'b00011_000110_00011;
        ingredient_text[11][0] = 16'b00011_000110_00011;
        ingredient_text[11][1] = 16'b00011_000110_00011;
        ingredient_text[11][2] = 16'b00011_000110_00011;
        ingredient_text[11][3] = 16'b00011_000110_00011;
        ingredient_text[11][4] = 16'b00011_000110_00011;
        ingredient_text[11][5] = 16'b00011_000110_00011;
        ingredient_text[11][6] = 16'b00011_000110_00011;
        ingredient_text[11][7] = 16'b00011_000110_00011;
        ingredient_text[11][8] = 16'b00011_000110_00011;
        ingredient_text[11][9] = 16'b00011_000110_00011;
        ingredient_text[11][10] = 16'b00011_000110_00011;
        ingredient_text[11][11] = 16'b00011_000110_00011;
        ingredient_text[11][12] = 16'b00011_000110_00011;
        ingredient_text[11][13] = 16'b00011_000110_00011;
        ingredient_text[11][14] = 16'b00011_000110_00011;
        ingredient_text[11][15] = 16'b00011_000110_00011;
        ingredient_text[11][16] = 16'b00011_000110_00011;
        ingredient_text[11][17] = 16'b00011_000110_00011;
        ingredient_text[11][18] = 16'b11111_111111_11111;
        ingredient_text[11][19] = 16'b01110_011110_01110;
        ingredient_text[11][20] = 16'b00011_000110_00011;
        ingredient_text[11][21] = 16'b00011_000110_00011;
        ingredient_text[11][22] = 16'b00011_000110_00011;
        ingredient_text[11][23] = 16'b00011_000110_00011;
        ingredient_text[11][24] = 16'b00011_000110_00011;
        ingredient_text[11][25] = 16'b00011_000110_00011;
        ingredient_text[11][26] = 16'b00011_000110_00011;
        ingredient_text[11][27] = 16'b00011_000110_00011;
        ingredient_text[11][28] = 16'b00011_000110_00011;
        ingredient_text[11][29] = 16'b00011_000110_00011;
        ingredient_text[11][30] = 16'b00011_000110_00011;
        ingredient_text[11][31] = 16'b00011_000110_00011;
        ingredient_text[11][32] = 16'b00011_000110_00011;
        ingredient_text[11][33] = 16'b00011_000110_00011;
        ingredient_text[11][34] = 16'b00011_000110_00011;
        ingredient_text[11][35] = 16'b00011_000110_00011;
        ingredient_text[11][36] = 16'b11111_111111_11111;
        ingredient_text[11][37] = 16'b11011_110111_11011;
        ingredient_text[11][38] = 16'b00011_000110_00011;
        ingredient_text[11][39] = 16'b11011_110111_11011;
        ingredient_text[11][40] = 16'b11111_111111_11111;
        ingredient_text[11][41] = 16'b00011_000110_00011;
        ingredient_text[11][42] = 16'b00011_000110_00011;
        ingredient_text[11][43] = 16'b00011_000110_00011;
        ingredient_text[11][44] = 16'b00011_000110_00011;
        ingredient_text[11][45] = 16'b00011_000110_00011;
        ingredient_text[11][46] = 16'b00011_000110_00011;
        ingredient_text[11][47] = 16'b00011_000110_00011;
        ingredient_text[11][48] = 16'b00011_000110_00011;
        ingredient_text[11][49] = 16'b00011_000110_00011;
        ingredient_text[11][50] = 16'b00011_000110_00011;
        ingredient_text[11][51] = 16'b00011_000110_00011;
        ingredient_text[11][52] = 16'b00011_000110_00011;
        ingredient_text[11][53] = 16'b00011_000110_00011;
        ingredient_text[11][54] = 16'b00011_000110_00011;
        ingredient_text[11][55] = 16'b00011_000110_00011;
        ingredient_text[11][56] = 16'b00011_000110_00011;
        ingredient_text[11][57] = 16'b00011_000110_00011;
        ingredient_text[11][58] = 16'b00011_000110_00011;
        ingredient_text[11][59] = 16'b00011_000110_00011;
        ingredient_text[11][60] = 16'b00011_000110_00011;
        ingredient_text[11][61] = 16'b00011_000110_00011;
        ingredient_text[11][62] = 16'b00011_000110_00011;
        ingredient_text[11][63] = 16'b00011_000110_00011;
        ingredient_text[11][64] = 16'b00011_000110_00011;
        ingredient_text[11][65] = 16'b00011_000110_00011;
        ingredient_text[11][66] = 16'b00011_000110_00011;
        ingredient_text[11][67] = 16'b00011_000110_00011;
        ingredient_text[11][68] = 16'b00011_000110_00011;
        ingredient_text[11][69] = 16'b00011_000110_00011;
        ingredient_text[11][70] = 16'b00011_000110_00011;
        ingredient_text[11][71] = 16'b00011_000110_00011;
        ingredient_text[11][72] = 16'b00011_000110_00011;
        ingredient_text[11][73] = 16'b11111_111111_11111;
        ingredient_text[11][74] = 16'b11111_111111_11111;
        ingredient_text[11][75] = 16'b00011_000110_00011;
        ingredient_text[11][76] = 16'b00011_000110_00011;
        ingredient_text[11][77] = 16'b00011_000110_00011;
        ingredient_text[11][78] = 16'b00011_000110_00011;
        ingredient_text[11][79] = 16'b00011_000110_00011;
        ingredient_text[12][0] = 16'b00011_000110_00011;
        ingredient_text[12][1] = 16'b00011_000110_00011;
        ingredient_text[12][2] = 16'b00011_000110_00011;
        ingredient_text[12][3] = 16'b00011_000110_00011;
        ingredient_text[12][4] = 16'b00011_000110_00011;
        ingredient_text[12][5] = 16'b00011_000110_00011;
        ingredient_text[12][6] = 16'b00011_000110_00011;
        ingredient_text[12][7] = 16'b00011_000110_00011;
        ingredient_text[12][8] = 16'b00011_000110_00011;
        ingredient_text[12][9] = 16'b00011_000110_00011;
        ingredient_text[12][10] = 16'b00011_000110_00011;
        ingredient_text[12][11] = 16'b00011_000110_00011;
        ingredient_text[12][12] = 16'b00011_000110_00011;
        ingredient_text[12][13] = 16'b00011_000110_00011;
        ingredient_text[12][14] = 16'b00011_000110_00011;
        ingredient_text[12][15] = 16'b00011_000110_00011;
        ingredient_text[12][16] = 16'b00011_000110_00011;
        ingredient_text[12][17] = 16'b00011_000110_00011;
        ingredient_text[12][18] = 16'b00011_000110_00011;
        ingredient_text[12][19] = 16'b00011_000110_00011;
        ingredient_text[12][20] = 16'b00011_000110_00011;
        ingredient_text[12][21] = 16'b00011_000110_00011;
        ingredient_text[12][22] = 16'b00011_000110_00011;
        ingredient_text[12][23] = 16'b00011_000110_00011;
        ingredient_text[12][24] = 16'b00011_000110_00011;
        ingredient_text[12][25] = 16'b00011_000110_00011;
        ingredient_text[12][26] = 16'b00011_000110_00011;
        ingredient_text[12][27] = 16'b00011_000110_00011;
        ingredient_text[12][28] = 16'b00011_000110_00011;
        ingredient_text[12][29] = 16'b00011_000110_00011;
        ingredient_text[12][30] = 16'b00011_000110_00011;
        ingredient_text[12][31] = 16'b00011_000110_00011;
        ingredient_text[12][32] = 16'b00011_000110_00011;
        ingredient_text[12][33] = 16'b00011_000110_00011;
        ingredient_text[12][34] = 16'b00011_000110_00011;
        ingredient_text[12][35] = 16'b00011_000110_00011;
        ingredient_text[12][36] = 16'b11111_111111_11111;
        ingredient_text[12][37] = 16'b11111_111111_11111;
        ingredient_text[12][38] = 16'b00011_000110_00011;
        ingredient_text[12][39] = 16'b11011_110111_11011;
        ingredient_text[12][40] = 16'b11111_111111_11111;
        ingredient_text[12][41] = 16'b00011_000110_00011;
        ingredient_text[12][42] = 16'b00011_000110_00011;
        ingredient_text[12][43] = 16'b00011_000110_00011;
        ingredient_text[12][44] = 16'b00011_000110_00011;
        ingredient_text[12][45] = 16'b00011_000110_00011;
        ingredient_text[12][46] = 16'b00011_000110_00011;
        ingredient_text[12][47] = 16'b00011_000110_00011;
        ingredient_text[12][48] = 16'b00011_000110_00011;
        ingredient_text[12][49] = 16'b00011_000110_00011;
        ingredient_text[12][50] = 16'b00011_000110_00011;
        ingredient_text[12][51] = 16'b00011_000110_00011;
        ingredient_text[12][52] = 16'b00011_000110_00011;
        ingredient_text[12][53] = 16'b00011_000110_00011;
        ingredient_text[12][54] = 16'b00011_000110_00011;
        ingredient_text[12][55] = 16'b00011_000110_00011;
        ingredient_text[12][56] = 16'b00011_000110_00011;
        ingredient_text[12][57] = 16'b00011_000110_00011;
        ingredient_text[12][58] = 16'b00011_000110_00011;
        ingredient_text[12][59] = 16'b00011_000110_00011;
        ingredient_text[12][60] = 16'b00011_000110_00011;
        ingredient_text[12][61] = 16'b00011_000110_00011;
        ingredient_text[12][62] = 16'b00011_000110_00011;
        ingredient_text[12][63] = 16'b00011_000110_00011;
        ingredient_text[12][64] = 16'b00011_000110_00011;
        ingredient_text[12][65] = 16'b00011_000110_00011;
        ingredient_text[12][66] = 16'b00011_000110_00011;
        ingredient_text[12][67] = 16'b00011_000110_00011;
        ingredient_text[12][68] = 16'b00011_000110_00011;
        ingredient_text[12][69] = 16'b00011_000110_00011;
        ingredient_text[12][70] = 16'b00011_000110_00011;
        ingredient_text[12][71] = 16'b00011_000110_00011;
        ingredient_text[12][72] = 16'b00011_000110_00011;
        ingredient_text[12][73] = 16'b11111_111111_11111;
        ingredient_text[12][74] = 16'b11011_110111_11011;
        ingredient_text[12][75] = 16'b00011_000110_00011;
        ingredient_text[12][76] = 16'b00011_000110_00011;
        ingredient_text[12][77] = 16'b00011_000110_00011;
        ingredient_text[12][78] = 16'b00011_000110_00011;
        ingredient_text[12][79] = 16'b00011_000110_00011;
        ingredient_text[13][0] = 16'b00011_000110_00011;
        ingredient_text[13][1] = 16'b00011_000110_00011;
        ingredient_text[13][2] = 16'b00011_000110_00011;
        ingredient_text[13][3] = 16'b00011_000110_00011;
        ingredient_text[13][4] = 16'b00011_000110_00011;
        ingredient_text[13][5] = 16'b00011_000110_00011;
        ingredient_text[13][6] = 16'b00011_000110_00011;
        ingredient_text[13][7] = 16'b00011_000110_00011;
        ingredient_text[13][8] = 16'b00011_000110_00011;
        ingredient_text[13][9] = 16'b00011_000110_00011;
        ingredient_text[13][10] = 16'b00011_000110_00011;
        ingredient_text[13][11] = 16'b00011_000110_00011;
        ingredient_text[13][12] = 16'b00011_000110_00011;
        ingredient_text[13][13] = 16'b00011_000110_00011;
        ingredient_text[13][14] = 16'b00011_000110_00011;
        ingredient_text[13][15] = 16'b00011_000110_00011;
        ingredient_text[13][16] = 16'b00011_000110_00011;
        ingredient_text[13][17] = 16'b00011_000110_00011;
        ingredient_text[13][18] = 16'b00011_000110_00011;
        ingredient_text[13][19] = 16'b00011_000110_00011;
        ingredient_text[13][20] = 16'b00011_000110_00011;
        ingredient_text[13][21] = 16'b00011_000110_00011;
        ingredient_text[13][22] = 16'b00011_000110_00011;
        ingredient_text[13][23] = 16'b00011_000110_00011;
        ingredient_text[13][24] = 16'b00011_000110_00011;
        ingredient_text[13][25] = 16'b00011_000110_00011;
        ingredient_text[13][26] = 16'b00011_000110_00011;
        ingredient_text[13][27] = 16'b00011_000110_00011;
        ingredient_text[13][28] = 16'b00011_000110_00011;
        ingredient_text[13][29] = 16'b00011_000110_00011;
        ingredient_text[13][30] = 16'b00011_000110_00011;
        ingredient_text[13][31] = 16'b00011_000110_00011;
        ingredient_text[13][32] = 16'b00011_000110_00011;
        ingredient_text[13][33] = 16'b00011_000110_00011;
        ingredient_text[13][34] = 16'b00011_000110_00011;
        ingredient_text[13][35] = 16'b00011_000110_00011;
        ingredient_text[13][36] = 16'b00011_000110_00011;
        ingredient_text[13][37] = 16'b00011_000110_00011;
        ingredient_text[13][38] = 16'b00011_000110_00011;
        ingredient_text[13][39] = 16'b00011_000110_00011;
        ingredient_text[13][40] = 16'b00011_000110_00011;
        ingredient_text[13][41] = 16'b00011_000110_00011;
        ingredient_text[13][42] = 16'b00011_000110_00011;
        ingredient_text[13][43] = 16'b00011_000110_00011;
        ingredient_text[13][44] = 16'b00011_000110_00011;
        ingredient_text[13][45] = 16'b00011_000110_00011;
        ingredient_text[13][46] = 16'b00011_000110_00011;
        ingredient_text[13][47] = 16'b00011_000110_00011;
        ingredient_text[13][48] = 16'b00011_000110_00011;
        ingredient_text[13][49] = 16'b00011_000110_00011;
        ingredient_text[13][50] = 16'b00011_000110_00011;
        ingredient_text[13][51] = 16'b00011_000110_00011;
        ingredient_text[13][52] = 16'b00011_000110_00011;
        ingredient_text[13][53] = 16'b00011_000110_00011;
        ingredient_text[13][54] = 16'b00011_000110_00011;
        ingredient_text[13][55] = 16'b00011_000110_00011;
        ingredient_text[13][56] = 16'b00011_000110_00011;
        ingredient_text[13][57] = 16'b00011_000110_00011;
        ingredient_text[13][58] = 16'b00011_000110_00011;
        ingredient_text[13][59] = 16'b00011_000110_00011;
        ingredient_text[13][60] = 16'b00011_000110_00011;
        ingredient_text[13][61] = 16'b00011_000110_00011;
        ingredient_text[13][62] = 16'b00011_000110_00011;
        ingredient_text[13][63] = 16'b00011_000110_00011;
        ingredient_text[13][64] = 16'b00011_000110_00011;
        ingredient_text[13][65] = 16'b00011_000110_00011;
        ingredient_text[13][66] = 16'b00011_000110_00011;
        ingredient_text[13][67] = 16'b00011_000110_00011;
        ingredient_text[13][68] = 16'b00011_000110_00011;
        ingredient_text[13][69] = 16'b00011_000110_00011;
        ingredient_text[13][70] = 16'b00011_000110_00011;
        ingredient_text[13][71] = 16'b00011_000110_00011;
        ingredient_text[13][72] = 16'b00011_000110_00011;
        ingredient_text[13][73] = 16'b00011_000110_00011;
        ingredient_text[13][74] = 16'b00011_000110_00011;
        ingredient_text[13][75] = 16'b00011_000110_00011;
        ingredient_text[13][76] = 16'b00011_000110_00011;
        ingredient_text[13][77] = 16'b00011_000110_00011;
        ingredient_text[13][78] = 16'b00011_000110_00011;
        ingredient_text[13][79] = 16'b00011_000110_00011;
        ingredient_text[14][0] = 16'b00011_000110_00011;
        ingredient_text[14][1] = 16'b00011_000110_00011;
        ingredient_text[14][2] = 16'b00011_000110_00011;
        ingredient_text[14][3] = 16'b00011_000110_00011;
        ingredient_text[14][4] = 16'b00011_000110_00011;
        ingredient_text[14][5] = 16'b00011_000110_00011;
        ingredient_text[14][6] = 16'b00011_000110_00011;
        ingredient_text[14][7] = 16'b00011_000110_00011;
        ingredient_text[14][8] = 16'b00011_000110_00011;
        ingredient_text[14][9] = 16'b00011_000110_00011;
        ingredient_text[14][10] = 16'b00011_000110_00011;
        ingredient_text[14][11] = 16'b00011_000110_00011;
        ingredient_text[14][12] = 16'b00011_000110_00011;
        ingredient_text[14][13] = 16'b00011_000110_00011;
        ingredient_text[14][14] = 16'b00011_000110_00011;
        ingredient_text[14][15] = 16'b00011_000110_00011;
        ingredient_text[14][16] = 16'b00011_000110_00011;
        ingredient_text[14][17] = 16'b00011_000110_00011;
        ingredient_text[14][18] = 16'b00011_000110_00011;
        ingredient_text[14][19] = 16'b00011_000110_00011;
        ingredient_text[14][20] = 16'b00011_000110_00011;
        ingredient_text[14][21] = 16'b00011_000110_00011;
        ingredient_text[14][22] = 16'b00011_000110_00011;
        ingredient_text[14][23] = 16'b00011_000110_00011;
        ingredient_text[14][24] = 16'b00011_000110_00011;
        ingredient_text[14][25] = 16'b00011_000110_00011;
        ingredient_text[14][26] = 16'b00011_000110_00011;
        ingredient_text[14][27] = 16'b00011_000110_00011;
        ingredient_text[14][28] = 16'b00011_000110_00011;
        ingredient_text[14][29] = 16'b00011_000110_00011;
        ingredient_text[14][30] = 16'b00011_000110_00011;
        ingredient_text[14][31] = 16'b00011_000110_00011;
        ingredient_text[14][32] = 16'b00011_000110_00011;
        ingredient_text[14][33] = 16'b00011_000110_00011;
        ingredient_text[14][34] = 16'b00011_000110_00011;
        ingredient_text[14][35] = 16'b00011_000110_00011;
        ingredient_text[14][36] = 16'b00011_000110_00011;
        ingredient_text[14][37] = 16'b00011_000110_00011;
        ingredient_text[14][38] = 16'b00011_000110_00011;
        ingredient_text[14][39] = 16'b00011_000110_00011;
        ingredient_text[14][40] = 16'b00011_000110_00011;
        ingredient_text[14][41] = 16'b00011_000110_00011;
        ingredient_text[14][42] = 16'b00011_000110_00011;
        ingredient_text[14][43] = 16'b00011_000110_00011;
        ingredient_text[14][44] = 16'b00011_000110_00011;
        ingredient_text[14][45] = 16'b00011_000110_00011;
        ingredient_text[14][46] = 16'b00011_000110_00011;
        ingredient_text[14][47] = 16'b00011_000110_00011;
        ingredient_text[14][48] = 16'b00011_000110_00011;
        ingredient_text[14][49] = 16'b00011_000110_00011;
        ingredient_text[14][50] = 16'b00011_000110_00011;
        ingredient_text[14][51] = 16'b00011_000110_00011;
        ingredient_text[14][52] = 16'b00011_000110_00011;
        ingredient_text[14][53] = 16'b00011_000110_00011;
        ingredient_text[14][54] = 16'b00011_000110_00011;
        ingredient_text[14][55] = 16'b00011_000110_00011;
        ingredient_text[14][56] = 16'b00011_000110_00011;
        ingredient_text[14][57] = 16'b00011_000110_00011;
        ingredient_text[14][58] = 16'b00011_000110_00011;
        ingredient_text[14][59] = 16'b00011_000110_00011;
        ingredient_text[14][60] = 16'b00011_000110_00011;
        ingredient_text[14][61] = 16'b00011_000110_00011;
        ingredient_text[14][62] = 16'b00011_000110_00011;
        ingredient_text[14][63] = 16'b00011_000110_00011;
        ingredient_text[14][64] = 16'b00011_000110_00011;
        ingredient_text[14][65] = 16'b00011_000110_00011;
        ingredient_text[14][66] = 16'b00011_000110_00011;
        ingredient_text[14][67] = 16'b00011_000110_00011;
        ingredient_text[14][68] = 16'b00011_000110_00011;
        ingredient_text[14][69] = 16'b00011_000110_00011;
        ingredient_text[14][70] = 16'b00011_000110_00011;
        ingredient_text[14][71] = 16'b00011_000110_00011;
        ingredient_text[14][72] = 16'b00011_000110_00011;
        ingredient_text[14][73] = 16'b00011_000110_00011;
        ingredient_text[14][74] = 16'b00011_000110_00011;
        ingredient_text[14][75] = 16'b00011_000110_00011;
        ingredient_text[14][76] = 16'b00011_000110_00011;
        ingredient_text[14][77] = 16'b00011_000110_00011;
        ingredient_text[14][78] = 16'b00011_000110_00011;
        ingredient_text[14][79] = 16'b00011_000110_00011;
        ingredient_text[15][0] = 16'b00011_000110_00011;
        ingredient_text[15][1] = 16'b00011_000110_00011;
        ingredient_text[15][2] = 16'b00011_000110_00011;
        ingredient_text[15][3] = 16'b00011_000110_00011;
        ingredient_text[15][4] = 16'b00011_000110_00011;
        ingredient_text[15][5] = 16'b00011_000110_00011;
        ingredient_text[15][6] = 16'b00011_000110_00011;
        ingredient_text[15][7] = 16'b00011_000110_00011;
        ingredient_text[15][8] = 16'b00011_000110_00011;
        ingredient_text[15][9] = 16'b00011_000110_00011;
        ingredient_text[15][10] = 16'b00011_000110_00011;
        ingredient_text[15][11] = 16'b00011_000110_00011;
        ingredient_text[15][12] = 16'b00011_000110_00011;
        ingredient_text[15][13] = 16'b00011_000110_00011;
        ingredient_text[15][14] = 16'b00011_000110_00011;
        ingredient_text[15][15] = 16'b00011_000110_00011;
        ingredient_text[15][16] = 16'b00011_000110_00011;
        ingredient_text[15][17] = 16'b00011_000110_00011;
        ingredient_text[15][18] = 16'b00011_000110_00011;
        ingredient_text[15][19] = 16'b00011_000110_00011;
        ingredient_text[15][20] = 16'b00011_000110_00011;
        ingredient_text[15][21] = 16'b00011_000110_00011;
        ingredient_text[15][22] = 16'b00011_000110_00011;
        ingredient_text[15][23] = 16'b00011_000110_00011;
        ingredient_text[15][24] = 16'b00011_000110_00011;
        ingredient_text[15][25] = 16'b00011_000110_00011;
        ingredient_text[15][26] = 16'b00011_000110_00011;
        ingredient_text[15][27] = 16'b00011_000110_00011;
        ingredient_text[15][28] = 16'b00011_000110_00011;
        ingredient_text[15][29] = 16'b00011_000110_00011;
        ingredient_text[15][30] = 16'b00011_000110_00011;
        ingredient_text[15][31] = 16'b00011_000110_00011;
        ingredient_text[15][32] = 16'b00011_000110_00011;
        ingredient_text[15][33] = 16'b00011_000110_00011;
        ingredient_text[15][34] = 16'b00011_000110_00011;
        ingredient_text[15][35] = 16'b00011_000110_00011;
        ingredient_text[15][36] = 16'b00011_000110_00011;
        ingredient_text[15][37] = 16'b00011_000110_00011;
        ingredient_text[15][38] = 16'b00011_000110_00011;
        ingredient_text[15][39] = 16'b00011_000110_00011;
        ingredient_text[15][40] = 16'b00011_000110_00011;
        ingredient_text[15][41] = 16'b00011_000110_00011;
        ingredient_text[15][42] = 16'b00011_000110_00011;
        ingredient_text[15][43] = 16'b00011_000110_00011;
        ingredient_text[15][44] = 16'b00011_000110_00011;
        ingredient_text[15][45] = 16'b00011_000110_00011;
        ingredient_text[15][46] = 16'b00011_000110_00011;
        ingredient_text[15][47] = 16'b00011_000110_00011;
        ingredient_text[15][48] = 16'b00011_000110_00011;
        ingredient_text[15][49] = 16'b00011_000110_00011;
        ingredient_text[15][50] = 16'b00011_000110_00011;
        ingredient_text[15][51] = 16'b00011_000110_00011;
        ingredient_text[15][52] = 16'b00011_000110_00011;
        ingredient_text[15][53] = 16'b00011_000110_00011;
        ingredient_text[15][54] = 16'b00011_000110_00011;
        ingredient_text[15][55] = 16'b00011_000110_00011;
        ingredient_text[15][56] = 16'b00011_000110_00011;
        ingredient_text[15][57] = 16'b00011_000110_00011;
        ingredient_text[15][58] = 16'b00011_000110_00011;
        ingredient_text[15][59] = 16'b00011_000110_00011;
        ingredient_text[15][60] = 16'b00011_000110_00011;
        ingredient_text[15][61] = 16'b00011_000110_00011;
        ingredient_text[15][62] = 16'b00011_000110_00011;
        ingredient_text[15][63] = 16'b00011_000110_00011;
        ingredient_text[15][64] = 16'b00011_000110_00011;
        ingredient_text[15][65] = 16'b00011_000110_00011;
        ingredient_text[15][66] = 16'b00011_000110_00011;
        ingredient_text[15][67] = 16'b00011_000110_00011;
        ingredient_text[15][68] = 16'b00011_000110_00011;
        ingredient_text[15][69] = 16'b00011_000110_00011;
        ingredient_text[15][70] = 16'b00011_000110_00011;
        ingredient_text[15][71] = 16'b00011_000110_00011;
        ingredient_text[15][72] = 16'b00011_000110_00011;
        ingredient_text[15][73] = 16'b00011_000110_00011;
        ingredient_text[15][74] = 16'b00011_000110_00011;
        ingredient_text[15][75] = 16'b00011_000110_00011;
        ingredient_text[15][76] = 16'b00011_000110_00011;
        ingredient_text[15][77] = 16'b00011_000110_00011;
        ingredient_text[15][78] = 16'b00011_000110_00011;
        ingredient_text[15][79] = 16'b00011_000110_00011;
        ingredient_text[16][0] = 16'b00011_000110_00011;
        ingredient_text[16][1] = 16'b00011_000110_00011;
        ingredient_text[16][2] = 16'b00011_000110_00011;
        ingredient_text[16][3] = 16'b00011_000110_00011;
        ingredient_text[16][4] = 16'b00011_000110_00011;
        ingredient_text[16][5] = 16'b00011_000110_00011;
        ingredient_text[16][6] = 16'b00011_000110_00011;
        ingredient_text[16][7] = 16'b00011_000110_00011;
        ingredient_text[16][8] = 16'b00011_000110_00011;
        ingredient_text[16][9] = 16'b00011_000110_00011;
        ingredient_text[16][10] = 16'b00011_000110_00011;
        ingredient_text[16][11] = 16'b00011_000110_00011;
        ingredient_text[16][12] = 16'b00011_000110_00011;
        ingredient_text[16][13] = 16'b00011_000110_00011;
        ingredient_text[16][14] = 16'b00011_000110_00011;
        ingredient_text[16][15] = 16'b00011_000110_00011;
        ingredient_text[16][16] = 16'b00011_000110_00011;
        ingredient_text[16][17] = 16'b00011_000110_00011;
        ingredient_text[16][18] = 16'b00011_000110_00011;
        ingredient_text[16][19] = 16'b00011_000110_00011;
        ingredient_text[16][20] = 16'b00011_000110_00011;
        ingredient_text[16][21] = 16'b00011_000110_00011;
        ingredient_text[16][22] = 16'b00011_000110_00011;
        ingredient_text[16][23] = 16'b00011_000110_00011;
        ingredient_text[16][24] = 16'b00011_000110_00011;
        ingredient_text[16][25] = 16'b00011_000110_00011;
        ingredient_text[16][26] = 16'b00011_000110_00011;
        ingredient_text[16][27] = 16'b00011_000110_00011;
        ingredient_text[16][28] = 16'b00011_000110_00011;
        ingredient_text[16][29] = 16'b00011_000110_00011;
        ingredient_text[16][30] = 16'b00011_000110_00011;
        ingredient_text[16][31] = 16'b00011_000110_00011;
        ingredient_text[16][32] = 16'b00011_000110_00011;
        ingredient_text[16][33] = 16'b00011_000110_00011;
        ingredient_text[16][34] = 16'b00011_000110_00011;
        ingredient_text[16][35] = 16'b00011_000110_00011;
        ingredient_text[16][36] = 16'b00011_000110_00011;
        ingredient_text[16][37] = 16'b00011_000110_00011;
        ingredient_text[16][38] = 16'b00011_000110_00011;
        ingredient_text[16][39] = 16'b00011_000110_00011;
        ingredient_text[16][40] = 16'b00011_000110_00011;
        ingredient_text[16][41] = 16'b00011_000110_00011;
        ingredient_text[16][42] = 16'b00011_000110_00011;
        ingredient_text[16][43] = 16'b00011_000110_00011;
        ingredient_text[16][44] = 16'b00011_000110_00011;
        ingredient_text[16][45] = 16'b00011_000110_00011;
        ingredient_text[16][46] = 16'b00011_000110_00011;
        ingredient_text[16][47] = 16'b00011_000110_00011;
        ingredient_text[16][48] = 16'b00011_000110_00011;
        ingredient_text[16][49] = 16'b00011_000110_00011;
        ingredient_text[16][50] = 16'b00011_000110_00011;
        ingredient_text[16][51] = 16'b00011_000110_00011;
        ingredient_text[16][52] = 16'b00011_000110_00011;
        ingredient_text[16][53] = 16'b00011_000110_00011;
        ingredient_text[16][54] = 16'b00011_000110_00011;
        ingredient_text[16][55] = 16'b00011_000110_00011;
        ingredient_text[16][56] = 16'b00011_000110_00011;
        ingredient_text[16][57] = 16'b00011_000110_00011;
        ingredient_text[16][58] = 16'b00011_000110_00011;
        ingredient_text[16][59] = 16'b00011_000110_00011;
        ingredient_text[16][60] = 16'b00011_000110_00011;
        ingredient_text[16][61] = 16'b00011_000110_00011;
        ingredient_text[16][62] = 16'b00011_000110_00011;
        ingredient_text[16][63] = 16'b00011_000110_00011;
        ingredient_text[16][64] = 16'b00011_000110_00011;
        ingredient_text[16][65] = 16'b00011_000110_00011;
        ingredient_text[16][66] = 16'b00011_000110_00011;
        ingredient_text[16][67] = 16'b00011_000110_00011;
        ingredient_text[16][68] = 16'b00011_000110_00011;
        ingredient_text[16][69] = 16'b00011_000110_00011;
        ingredient_text[16][70] = 16'b00011_000110_00011;
        ingredient_text[16][71] = 16'b00011_000110_00011;
        ingredient_text[16][72] = 16'b00011_000110_00011;
        ingredient_text[16][73] = 16'b00011_000110_00011;
        ingredient_text[16][74] = 16'b00011_000110_00011;
        ingredient_text[16][75] = 16'b00011_000110_00011;
        ingredient_text[16][76] = 16'b00011_000110_00011;
        ingredient_text[16][77] = 16'b00011_000110_00011;
        ingredient_text[16][78] = 16'b00011_000110_00011;
        ingredient_text[16][79] = 16'b00011_000110_00011;



        
        //ingredient
        rice_raw[0][0] = 16'b11111_111110_11111;
        rice_raw[0][1] = 16'b11111_111110_11111;
        rice_raw[0][2] = 16'b11111_111110_11111;
        rice_raw[0][3] = 16'b11111_111110_11111;
        rice_raw[0][4] = 16'b11111_111110_11111;
        rice_raw[0][5] = 16'b11111_111110_11111;
        rice_raw[0][6] = 16'b11111_111110_11111;
        rice_raw[0][7] = 16'b11111_111110_11111;
        rice_raw[0][8] = 16'b11111_111110_11111;
        rice_raw[0][9] = 16'b11111_111110_11111;
        rice_raw[0][10] = 16'b11111_111110_11111;
        rice_raw[0][11] = 16'b11111_111110_11111;
        rice_raw[0][12] = 16'b11111_111110_11111;
        rice_raw[0][13] = 16'b11111_111110_11111;
        rice_raw[0][14] = 16'b11111_111110_11111;
        rice_raw[1][0] = 16'b11111_111110_11111;
        rice_raw[1][1] = 16'b00000_000000_00000;
        rice_raw[1][2] = 16'b00000_000000_00000;
        rice_raw[1][3] = 16'b00000_000000_00000;
        rice_raw[1][4] = 16'b00000_000000_00000;
        rice_raw[1][5] = 16'b00000_000000_00000;
        rice_raw[1][6] = 16'b00000_000000_00000;
        rice_raw[1][7] = 16'b00000_000000_00000;
        rice_raw[1][8] = 16'b00000_000000_00000;
        rice_raw[1][9] = 16'b00000_000000_00000;
        rice_raw[1][10] = 16'b00000_000000_00000;
        rice_raw[1][11] = 16'b00000_000000_00000;
        rice_raw[1][12] = 16'b00000_000000_00000;
        rice_raw[1][13] = 16'b00000_000000_00000;
        rice_raw[1][14] = 16'b11111_111110_11111;
        rice_raw[2][0] = 16'b11111_111110_11111;
        rice_raw[2][1] = 16'b00000_000000_00000;
        rice_raw[2][2] = 16'b00000_000000_00000;
        rice_raw[2][3] = 16'b00000_000000_00000;
        rice_raw[2][4] = 16'b00000_000000_00000;
        rice_raw[2][5] = 16'b00000_000000_00000;
        rice_raw[2][6] = 16'b00000_110000_11111;
        rice_raw[2][7] = 16'b00000_110000_11111;
        rice_raw[2][8] = 16'b00000_110000_11111;
        rice_raw[2][9] = 16'b00000_000000_00000;
        rice_raw[2][10] = 16'b00000_000000_00000;
        rice_raw[2][11] = 16'b00000_000000_00000;
        rice_raw[2][12] = 16'b00000_000000_00000;
        rice_raw[2][13] = 16'b00000_000000_00000;
        rice_raw[2][14] = 16'b11111_111110_11111;
        rice_raw[3][0] = 16'b11111_111110_11111;
        rice_raw[3][1] = 16'b00000_000000_00000;
        rice_raw[3][2] = 16'b00000_000000_00000;
        rice_raw[3][3] = 16'b00000_110000_11111;
        rice_raw[3][4] = 16'b00000_110000_11111;
        rice_raw[3][5] = 16'b00000_110000_11111;
        rice_raw[3][6] = 16'b00000_110000_11111;
        rice_raw[3][7] = 16'b00000_110000_11111;
        rice_raw[3][8] = 16'b00000_110000_11111;
        rice_raw[3][9] = 16'b00000_110000_11111;
        rice_raw[3][10] = 16'b00000_110000_11111;
        rice_raw[3][11] = 16'b00000_110000_11111;
        rice_raw[3][12] = 16'b00000_000000_00000;
        rice_raw[3][13] = 16'b00000_000000_00000;
        rice_raw[3][14] = 16'b11111_111110_11111;
        rice_raw[4][0] = 16'b11111_111110_11111;
        rice_raw[4][1] = 16'b00000_000000_00000;
        rice_raw[4][2] = 16'b00000_000000_00000;
        rice_raw[4][3] = 16'b00000_110000_11111;
        rice_raw[4][4] = 16'b00000_110000_11111;
        rice_raw[4][5] = 16'b00000_110000_11111;
        rice_raw[4][6] = 16'b00000_110000_11111;
        rice_raw[4][7] = 16'b00000_110000_11111;
        rice_raw[4][8] = 16'b00000_110000_11111;
        rice_raw[4][9] = 16'b00000_110000_11111;
        rice_raw[4][10] = 16'b00000_110000_11111;
        rice_raw[4][11] = 16'b00000_110000_11111;
        rice_raw[4][12] = 16'b00000_000000_00000;
        rice_raw[4][13] = 16'b00000_000000_00000;
        rice_raw[4][14] = 16'b11111_111110_11111;
        rice_raw[5][0] = 16'b11111_111110_11111;
        rice_raw[5][1] = 16'b00000_000000_00000;
        rice_raw[5][2] = 16'b00000_110000_11111;
        rice_raw[5][3] = 16'b00000_110000_11111;
        rice_raw[5][4] = 16'b00000_110000_11111;
        rice_raw[5][5] = 16'b00000_110000_11111;
        rice_raw[5][6] = 16'b00000_110000_11111;
        rice_raw[5][7] = 16'b00000_110000_11111;
        rice_raw[5][8] = 16'b00000_110000_11111;
        rice_raw[5][9] = 16'b00000_110000_11111;
        rice_raw[5][10] = 16'b00000_110000_11111;
        rice_raw[5][11] = 16'b00000_110000_11111;
        rice_raw[5][12] = 16'b00000_110000_11111;
        rice_raw[5][13] = 16'b00000_000000_00000;
        rice_raw[5][14] = 16'b11111_111110_11111;
        rice_raw[6][0] = 16'b11111_111110_11111;
        rice_raw[6][1] = 16'b00000_000000_00000;
        rice_raw[6][2] = 16'b00000_110000_11111;
        rice_raw[6][3] = 16'b00000_110000_11111;
        rice_raw[6][4] = 16'b11111_111110_11111;
        rice_raw[6][5] = 16'b11111_111110_11111;
        rice_raw[6][6] = 16'b10001_100011_10001;
        rice_raw[6][7] = 16'b11111_111110_11111;
        rice_raw[6][8] = 16'b11111_111110_11111;
        rice_raw[6][9] = 16'b11111_111110_11111;
        rice_raw[6][10] = 16'b11111_111110_11111;
        rice_raw[6][11] = 16'b00000_110000_11111;
        rice_raw[6][12] = 16'b00000_110000_11111;
        rice_raw[6][13] = 16'b00000_000000_00000;
        rice_raw[6][14] = 16'b11111_111110_11111;
        rice_raw[7][0] = 16'b11111_111110_11111;
        rice_raw[7][1] = 16'b00000_000000_00000;
        rice_raw[7][2] = 16'b00000_110000_11111;
        rice_raw[7][3] = 16'b11111_111110_11111;
        rice_raw[7][4] = 16'b11111_111110_11111;
        rice_raw[7][5] = 16'b11111_111110_11111;
        rice_raw[7][6] = 16'b11111_111110_11111;
        rice_raw[7][7] = 16'b11111_111110_11111;
        rice_raw[7][8] = 16'b11111_111110_11111;
        rice_raw[7][9] = 16'b10001_100011_10001;
        rice_raw[7][10] = 16'b11111_111110_11111;
        rice_raw[7][11] = 16'b11111_111110_11111;
        rice_raw[7][12] = 16'b00000_110000_11111;
        rice_raw[7][13] = 16'b00000_000000_00000;
        rice_raw[7][14] = 16'b11111_111110_11111;
        rice_raw[8][0] = 16'b11111_111110_11111;
        rice_raw[8][1] = 16'b00000_000000_00000;
        rice_raw[8][2] = 16'b00000_000000_00000;
        rice_raw[8][3] = 16'b10001_100011_10001;
        rice_raw[8][4] = 16'b11111_111110_11111;
        rice_raw[8][5] = 16'b10001_100011_10001;
        rice_raw[8][6] = 16'b11111_111110_11111;
        rice_raw[8][7] = 16'b10001_100011_10001;
        rice_raw[8][8] = 16'b11111_111110_11111;
        rice_raw[8][9] = 16'b11111_111110_11111;
        rice_raw[8][10] = 16'b11111_111110_11111;
        rice_raw[8][11] = 16'b10001_100011_10001;
        rice_raw[8][12] = 16'b00000_000000_00000;
        rice_raw[8][13] = 16'b00000_000000_00000;
        rice_raw[8][14] = 16'b11111_111110_11111;
        rice_raw[9][0] = 16'b11111_111110_11111;
        rice_raw[9][1] = 16'b00000_000000_00000;
        rice_raw[9][2] = 16'b00000_000000_00000;
        rice_raw[9][3] = 16'b11111_111110_11111;
        rice_raw[9][4] = 16'b11111_111110_11111;
        rice_raw[9][5] = 16'b11111_111110_11111;
        rice_raw[9][6] = 16'b11111_111110_11111;
        rice_raw[9][7] = 16'b11111_111110_11111;
        rice_raw[9][8] = 16'b11111_111110_11111;
        rice_raw[9][9] = 16'b10001_100011_10001;
        rice_raw[9][10] = 16'b11111_111110_11111;
        rice_raw[9][11] = 16'b11111_111110_11111;
        rice_raw[9][12] = 16'b00000_000000_00000;
        rice_raw[9][13] = 16'b00000_000000_00000;
        rice_raw[9][14] = 16'b11111_111110_11111;
        rice_raw[10][0] = 16'b11111_111110_11111;
        rice_raw[10][1] = 16'b00000_000000_00000;
        rice_raw[10][2] = 16'b00000_000000_00000;
        rice_raw[10][3] = 16'b00000_000000_00000;
        rice_raw[10][4] = 16'b11111_111110_11111;
        rice_raw[10][5] = 16'b11111_111110_11111;
        rice_raw[10][6] = 16'b10001_100011_10001;
        rice_raw[10][7] = 16'b11111_111110_11111;
        rice_raw[10][8] = 16'b11111_111110_11111;
        rice_raw[10][9] = 16'b11111_111110_11111;
        rice_raw[10][10] = 16'b11111_111110_11111;
        rice_raw[10][11] = 16'b00000_000000_00000;
        rice_raw[10][12] = 16'b00000_000000_00000;
        rice_raw[10][13] = 16'b00000_000000_00000;
        rice_raw[10][14] = 16'b11111_111110_11111;
        rice_raw[11][0] = 16'b11111_111110_11111;
        rice_raw[11][1] = 16'b00000_000000_00000;
        rice_raw[11][2] = 16'b00000_000000_00000;
        rice_raw[11][3] = 16'b00000_000000_00000;
        rice_raw[11][4] = 16'b00000_000000_00000;
        rice_raw[11][5] = 16'b11111_111110_11111;
        rice_raw[11][6] = 16'b11111_111110_11111;
        rice_raw[11][7] = 16'b11111_111110_11111;
        rice_raw[11][8] = 16'b10001_100011_10001;
        rice_raw[11][9] = 16'b11111_111110_11111;
        rice_raw[11][10] = 16'b00000_000000_00000;
        rice_raw[11][11] = 16'b00000_000000_00000;
        rice_raw[11][12] = 16'b00000_000000_00000;
        rice_raw[11][13] = 16'b00000_000000_00000;
        rice_raw[11][14] = 16'b11111_111110_11111;
        rice_raw[12][0] = 16'b11111_111110_11111;
        rice_raw[12][1] = 16'b00000_000000_00000;
        rice_raw[12][2] = 16'b00000_000000_00000;
        rice_raw[12][3] = 16'b00000_000000_00000;
        rice_raw[12][4] = 16'b00000_000000_00000;
        rice_raw[12][5] = 16'b00000_000000_00000;
        rice_raw[12][6] = 16'b11111_111110_11111;
        rice_raw[12][7] = 16'b11111_111110_11111;
        rice_raw[12][8] = 16'b11111_111110_11111;
        rice_raw[12][9] = 16'b00000_000000_00000;
        rice_raw[12][10] = 16'b00000_000000_00000;
        rice_raw[12][11] = 16'b00000_000000_00000;
        rice_raw[12][12] = 16'b00000_000000_00000;
        rice_raw[12][13] = 16'b00000_000000_00000;
        rice_raw[12][14] = 16'b11111_111110_11111;
        rice_raw[13][0] = 16'b11111_111110_11111;
        rice_raw[13][1] = 16'b00000_000000_00000;
        rice_raw[13][2] = 16'b00000_000000_00000;
        rice_raw[13][3] = 16'b00000_000000_00000;
        rice_raw[13][4] = 16'b00000_000000_00000;
        rice_raw[13][5] = 16'b00000_000000_00000;
        rice_raw[13][6] = 16'b00000_000000_00000;
        rice_raw[13][7] = 16'b00000_000000_00000;
        rice_raw[13][8] = 16'b00000_000000_00000;
        rice_raw[13][9] = 16'b00000_000000_00000;
        rice_raw[13][10] = 16'b00000_000000_00000;
        rice_raw[13][11] = 16'b00000_000000_00000;
        rice_raw[13][12] = 16'b00000_000000_00000;
        rice_raw[13][13] = 16'b00000_000000_00000;
        rice_raw[13][14] = 16'b11111_111110_11111;
        rice_raw[14][0] = 16'b11111_111110_11111;
        rice_raw[14][1] = 16'b11111_111110_11111;
        rice_raw[14][2] = 16'b11111_111110_11111;
        rice_raw[14][3] = 16'b11111_111110_11111;
        rice_raw[14][4] = 16'b11111_111110_11111;
        rice_raw[14][5] = 16'b11111_111110_11111;
        rice_raw[14][6] = 16'b11111_111110_11111;
        rice_raw[14][7] = 16'b11111_111110_11111;
        rice_raw[14][8] = 16'b11111_111110_11111;
        rice_raw[14][9] = 16'b11111_111110_11111;
        rice_raw[14][10] = 16'b11111_111110_11111;
        rice_raw[14][11] = 16'b11111_111110_11111;
        rice_raw[14][12] = 16'b11111_111110_11111;
        rice_raw[14][13] = 16'b11111_111110_11111;
        rice_raw[14][14] = 16'b11111_111110_11111;

        
        rice_boiled[0][0] = 16'b00000_000110_11111;
        rice_boiled[0][1] = 16'b00000_000110_11111;
        rice_boiled[0][2] = 16'b00000_000110_11111;
        rice_boiled[0][3] = 16'b00000_000110_11111;
        rice_boiled[0][4] = 16'b00000_000110_11111;
        rice_boiled[0][5] = 16'b00000_000110_11111;
        rice_boiled[0][6] = 16'b00000_000110_11111;
        rice_boiled[0][7] = 16'b00000_000110_11111;
        rice_boiled[0][8] = 16'b00000_000110_11111;
        rice_boiled[0][9] = 16'b00000_000110_11111;
        rice_boiled[0][10] = 16'b00000_000110_11111;
        rice_boiled[0][11] = 16'b00000_000110_11111;
        rice_boiled[0][12] = 16'b00000_000110_11111;
        rice_boiled[0][13] = 16'b00000_000110_11111;
        rice_boiled[0][14] = 16'b00000_000110_11111;
        rice_boiled[1][0] = 16'b00000_000110_11111;
        rice_boiled[1][1] = 16'b00000_000000_00000;
        rice_boiled[1][2] = 16'b00000_000000_00000;
        rice_boiled[1][3] = 16'b00000_000000_00000;
        rice_boiled[1][4] = 16'b00000_000000_00000;
        rice_boiled[1][5] = 16'b00000_000000_00000;
        rice_boiled[1][6] = 16'b00000_000000_00000;
        rice_boiled[1][7] = 16'b00000_000000_00000;
        rice_boiled[1][8] = 16'b00000_000000_00000;
        rice_boiled[1][9] = 16'b00000_000000_00000;
        rice_boiled[1][10] = 16'b00000_000000_00000;
        rice_boiled[1][11] = 16'b00000_000000_00000;
        rice_boiled[1][12] = 16'b00000_000000_00000;
        rice_boiled[1][13] = 16'b00000_000000_00000;
        rice_boiled[1][14] = 16'b00000_000110_11111;
        rice_boiled[2][0] = 16'b00000_000110_11111;
        rice_boiled[2][1] = 16'b00000_000000_00000;
        rice_boiled[2][2] = 16'b00000_000000_00000;
        rice_boiled[2][3] = 16'b00000_000000_00000;
        rice_boiled[2][4] = 16'b00000_000000_00000;
        rice_boiled[2][5] = 16'b00000_000000_00000;
        rice_boiled[2][6] = 16'b00000_110000_11111;
        rice_boiled[2][7] = 16'b00000_110000_11111;
        rice_boiled[2][8] = 16'b00000_110000_11111;
        rice_boiled[2][9] = 16'b00000_000000_00000;
        rice_boiled[2][10] = 16'b00000_000000_00000;
        rice_boiled[2][11] = 16'b00000_000000_00000;
        rice_boiled[2][12] = 16'b00000_000000_00000;
        rice_boiled[2][13] = 16'b00000_000000_00000;
        rice_boiled[2][14] = 16'b00000_000110_11111;
        rice_boiled[3][0] = 16'b00000_000110_11111;
        rice_boiled[3][1] = 16'b00000_000000_00000;
        rice_boiled[3][2] = 16'b00000_000000_00000;
        rice_boiled[3][3] = 16'b00000_110000_11111;
        rice_boiled[3][4] = 16'b00000_110000_11111;
        rice_boiled[3][5] = 16'b00000_110000_11111;
        rice_boiled[3][6] = 16'b00000_110000_11111;
        rice_boiled[3][7] = 16'b00000_110000_11111;
        rice_boiled[3][8] = 16'b00000_110000_11111;
        rice_boiled[3][9] = 16'b00000_110000_11111;
        rice_boiled[3][10] = 16'b00000_110000_11111;
        rice_boiled[3][11] = 16'b00000_110000_11111;
        rice_boiled[3][12] = 16'b00000_000000_00000;
        rice_boiled[3][13] = 16'b00000_000000_00000;
        rice_boiled[3][14] = 16'b00000_000110_11111;
        rice_boiled[4][0] = 16'b00000_000110_11111;
        rice_boiled[4][1] = 16'b00000_000000_00000;
        rice_boiled[4][2] = 16'b00000_000000_00000;
        rice_boiled[4][3] = 16'b00000_110000_11111;
        rice_boiled[4][4] = 16'b00000_110000_11111;
        rice_boiled[4][5] = 16'b00000_110000_11111;
        rice_boiled[4][6] = 16'b00000_110000_11111;
        rice_boiled[4][7] = 16'b00000_110000_11111;
        rice_boiled[4][8] = 16'b00000_110000_11111;
        rice_boiled[4][9] = 16'b00000_110000_11111;
        rice_boiled[4][10] = 16'b00000_110000_11111;
        rice_boiled[4][11] = 16'b00000_110000_11111;
        rice_boiled[4][12] = 16'b00000_000000_00000;
        rice_boiled[4][13] = 16'b00000_000000_00000;
        rice_boiled[4][14] = 16'b00000_000110_11111;
        rice_boiled[5][0] = 16'b00000_000110_11111;
        rice_boiled[5][1] = 16'b00000_000000_00000;
        rice_boiled[5][2] = 16'b00000_110000_11111;
        rice_boiled[5][3] = 16'b00000_110000_11111;
        rice_boiled[5][4] = 16'b00000_110000_11111;
        rice_boiled[5][5] = 16'b00000_110000_11111;
        rice_boiled[5][6] = 16'b00000_110000_11111;
        rice_boiled[5][7] = 16'b00000_110000_11111;
        rice_boiled[5][8] = 16'b00000_110000_11111;
        rice_boiled[5][9] = 16'b00000_110000_11111;
        rice_boiled[5][10] = 16'b00000_110000_11111;
        rice_boiled[5][11] = 16'b00000_110000_11111;
        rice_boiled[5][12] = 16'b00000_110000_11111;
        rice_boiled[5][13] = 16'b00000_000000_00000;
        rice_boiled[5][14] = 16'b00000_000110_11111;
        rice_boiled[6][0] = 16'b00000_000110_11111;
        rice_boiled[6][1] = 16'b00000_000000_00000;
        rice_boiled[6][2] = 16'b00000_110000_11111;
        rice_boiled[6][3] = 16'b00000_110000_11111;
        rice_boiled[6][4] = 16'b11111_111110_11111;
        rice_boiled[6][5] = 16'b11111_111110_11111;
        rice_boiled[6][6] = 16'b10001_100011_10001;
        rice_boiled[6][7] = 16'b11111_111110_11111;
        rice_boiled[6][8] = 16'b11111_111110_11111;
        rice_boiled[6][9] = 16'b11111_111110_11111;
        rice_boiled[6][10] = 16'b11111_111110_11111;
        rice_boiled[6][11] = 16'b00000_110000_11111;
        rice_boiled[6][12] = 16'b00000_110000_11111;
        rice_boiled[6][13] = 16'b00000_000000_00000;
        rice_boiled[6][14] = 16'b00000_000110_11111;
        rice_boiled[7][0] = 16'b00000_000110_11111;
        rice_boiled[7][1] = 16'b00000_000000_00000;
        rice_boiled[7][2] = 16'b00000_110000_11111;
        rice_boiled[7][3] = 16'b11111_111110_11111;
        rice_boiled[7][4] = 16'b11111_111110_11111;
        rice_boiled[7][5] = 16'b11111_111110_11111;
        rice_boiled[7][6] = 16'b11111_111110_11111;
        rice_boiled[7][7] = 16'b11111_111110_11111;
        rice_boiled[7][8] = 16'b11111_111110_11111;
        rice_boiled[7][9] = 16'b10001_100011_10001;
        rice_boiled[7][10] = 16'b11111_111110_11111;
        rice_boiled[7][11] = 16'b11111_111110_11111;
        rice_boiled[7][12] = 16'b00000_110000_11111;
        rice_boiled[7][13] = 16'b00000_000000_00000;
        rice_boiled[7][14] = 16'b00000_000110_11111;
        rice_boiled[8][0] = 16'b00000_000110_11111;
        rice_boiled[8][1] = 16'b00000_000000_00000;
        rice_boiled[8][2] = 16'b00000_000000_00000;
        rice_boiled[8][3] = 16'b10001_100011_10001;
        rice_boiled[8][4] = 16'b11111_111110_11111;
        rice_boiled[8][5] = 16'b10001_100011_10001;
        rice_boiled[8][6] = 16'b11111_111110_11111;
        rice_boiled[8][7] = 16'b10001_100011_10001;
        rice_boiled[8][8] = 16'b11111_111110_11111;
        rice_boiled[8][9] = 16'b11111_111110_11111;
        rice_boiled[8][10] = 16'b11111_111110_11111;
        rice_boiled[8][11] = 16'b10001_100011_10001;
        rice_boiled[8][12] = 16'b00000_000000_00000;
        rice_boiled[8][13] = 16'b00000_000000_00000;
        rice_boiled[8][14] = 16'b00000_000110_11111;
        rice_boiled[9][0] = 16'b00000_000110_11111;
        rice_boiled[9][1] = 16'b00000_000000_00000;
        rice_boiled[9][2] = 16'b00000_000000_00000;
        rice_boiled[9][3] = 16'b11111_111110_11111;
        rice_boiled[9][4] = 16'b11111_111110_11111;
        rice_boiled[9][5] = 16'b11111_111110_11111;
        rice_boiled[9][6] = 16'b11111_111110_11111;
        rice_boiled[9][7] = 16'b11111_111110_11111;
        rice_boiled[9][8] = 16'b11111_111110_11111;
        rice_boiled[9][9] = 16'b10001_100011_10001;
        rice_boiled[9][10] = 16'b11111_111110_11111;
        rice_boiled[9][11] = 16'b11111_111110_11111;
        rice_boiled[9][12] = 16'b00000_000000_00000;
        rice_boiled[9][13] = 16'b00000_000000_00000;
        rice_boiled[9][14] = 16'b00000_000110_11111;
        rice_boiled[10][0] = 16'b00000_000110_11111;
        rice_boiled[10][1] = 16'b00000_000000_00000;
        rice_boiled[10][2] = 16'b00000_000000_00000;
        rice_boiled[10][3] = 16'b00000_000000_00000;
        rice_boiled[10][4] = 16'b11111_111110_11111;
        rice_boiled[10][5] = 16'b11111_111110_11111;
        rice_boiled[10][6] = 16'b10001_100011_10001;
        rice_boiled[10][7] = 16'b11111_111110_11111;
        rice_boiled[10][8] = 16'b11111_111110_11111;
        rice_boiled[10][9] = 16'b11111_111110_11111;
        rice_boiled[10][10] = 16'b11111_111110_11111;
        rice_boiled[10][11] = 16'b00000_000000_00000;
        rice_boiled[10][12] = 16'b00000_000000_00000;
        rice_boiled[10][13] = 16'b00000_000000_00000;
        rice_boiled[10][14] = 16'b00000_000110_11111;
        rice_boiled[11][0] = 16'b00000_000110_11111;
        rice_boiled[11][1] = 16'b00000_000000_00000;
        rice_boiled[11][2] = 16'b00000_000000_00000;
        rice_boiled[11][3] = 16'b00000_000000_00000;
        rice_boiled[11][4] = 16'b00000_000000_00000;
        rice_boiled[11][5] = 16'b11111_111110_11111;
        rice_boiled[11][6] = 16'b11111_111110_11111;
        rice_boiled[11][7] = 16'b11111_111110_11111;
        rice_boiled[11][8] = 16'b10001_100011_10001;
        rice_boiled[11][9] = 16'b11111_111110_11111;
        rice_boiled[11][10] = 16'b00000_000000_00000;
        rice_boiled[11][11] = 16'b00000_000000_00000;
        rice_boiled[11][12] = 16'b00000_000000_00000;
        rice_boiled[11][13] = 16'b00000_000000_00000;
        rice_boiled[11][14] = 16'b00000_000110_11111;
        rice_boiled[12][0] = 16'b00000_000110_11111;
        rice_boiled[12][1] = 16'b00000_000000_00000;
        rice_boiled[12][2] = 16'b00000_000000_00000;
        rice_boiled[12][3] = 16'b00000_000000_00000;
        rice_boiled[12][4] = 16'b00000_000000_00000;
        rice_boiled[12][5] = 16'b00000_000000_00000;
        rice_boiled[12][6] = 16'b11111_111110_11111;
        rice_boiled[12][7] = 16'b11111_111110_11111;
        rice_boiled[12][8] = 16'b11111_111110_11111;
        rice_boiled[12][9] = 16'b00000_000000_00000;
        rice_boiled[12][10] = 16'b00000_000000_00000;
        rice_boiled[12][11] = 16'b00000_000000_00000;
        rice_boiled[12][12] = 16'b00000_000000_00000;
        rice_boiled[12][13] = 16'b00000_000000_00000;
        rice_boiled[12][14] = 16'b00000_000110_11111;
        rice_boiled[13][0] = 16'b00000_000110_11111;
        rice_boiled[13][1] = 16'b00000_000000_00000;
        rice_boiled[13][2] = 16'b00000_000000_00000;
        rice_boiled[13][3] = 16'b00000_000000_00000;
        rice_boiled[13][4] = 16'b00000_000000_00000;
        rice_boiled[13][5] = 16'b00000_000000_00000;
        rice_boiled[13][6] = 16'b00000_000000_00000;
        rice_boiled[13][7] = 16'b00000_000000_00000;
        rice_boiled[13][8] = 16'b00000_000000_00000;
        rice_boiled[13][9] = 16'b00000_000000_00000;
        rice_boiled[13][10] = 16'b00000_000000_00000;
        rice_boiled[13][11] = 16'b00000_000000_00000;
        rice_boiled[13][12] = 16'b00000_000000_00000;
        rice_boiled[13][13] = 16'b00000_000000_00000;
        rice_boiled[13][14] = 16'b00000_000110_11111;
        rice_boiled[14][0] = 16'b00000_000110_11111;
        rice_boiled[14][1] = 16'b00000_000110_11111;
        rice_boiled[14][2] = 16'b00000_000110_11111;
        rice_boiled[14][3] = 16'b00000_000110_11111;
        rice_boiled[14][4] = 16'b00000_000110_11111;
        rice_boiled[14][5] = 16'b00000_000110_11111;
        rice_boiled[14][6] = 16'b00000_000110_11111;
        rice_boiled[14][7] = 16'b00000_000110_11111;
        rice_boiled[14][8] = 16'b00000_000110_11111;
        rice_boiled[14][9] = 16'b00000_000110_11111;
        rice_boiled[14][10] = 16'b00000_000110_11111;
        rice_boiled[14][11] = 16'b00000_000110_11111;
        rice_boiled[14][12] = 16'b00000_000110_11111;
        rice_boiled[14][13] = 16'b00000_000110_11111;
        rice_boiled[14][14] = 16'b00000_000110_11111;

        
        rice_chopped[0][0] = 16'b00000_111111_00001;
        rice_chopped[0][1] = 16'b00000_111111_00001;
        rice_chopped[0][2] = 16'b00000_111111_00001;
        rice_chopped[0][3] = 16'b00000_111111_00001;
        rice_chopped[0][4] = 16'b00000_111111_00001;
        rice_chopped[0][5] = 16'b00000_111111_00001;
        rice_chopped[0][6] = 16'b00000_111111_00001;
        rice_chopped[0][7] = 16'b00000_111111_00001;
        rice_chopped[0][8] = 16'b00000_111111_00001;
        rice_chopped[0][9] = 16'b00000_111111_00001;
        rice_chopped[0][10] = 16'b00000_111111_00001;
        rice_chopped[0][11] = 16'b00000_111111_00001;
        rice_chopped[0][12] = 16'b00000_111111_00001;
        rice_chopped[0][13] = 16'b00000_111111_00001;
        rice_chopped[0][14] = 16'b00000_111111_00001;
        rice_chopped[1][0] = 16'b00000_111111_00001;
        rice_chopped[1][1] = 16'b00000_000000_00000;
        rice_chopped[1][2] = 16'b00000_000000_00000;
        rice_chopped[1][3] = 16'b00000_000000_00000;
        rice_chopped[1][4] = 16'b00000_000000_00000;
        rice_chopped[1][5] = 16'b00000_000000_00000;
        rice_chopped[1][6] = 16'b00000_000000_00000;
        rice_chopped[1][7] = 16'b00000_000000_00000;
        rice_chopped[1][8] = 16'b00000_000000_00000;
        rice_chopped[1][9] = 16'b00000_000000_00000;
        rice_chopped[1][10] = 16'b00000_000000_00000;
        rice_chopped[1][11] = 16'b00000_000000_00000;
        rice_chopped[1][12] = 16'b00000_000000_00000;
        rice_chopped[1][13] = 16'b00000_000000_00000;
        rice_chopped[1][14] = 16'b00000_111111_00001;
        rice_chopped[2][0] = 16'b00000_111111_00001;
        rice_chopped[2][1] = 16'b00000_000000_00000;
        rice_chopped[2][2] = 16'b00000_000000_00000;
        rice_chopped[2][3] = 16'b00000_000000_00000;
        rice_chopped[2][4] = 16'b00000_000000_00000;
        rice_chopped[2][5] = 16'b00000_000000_00000;
        rice_chopped[2][6] = 16'b00000_110000_11111;
        rice_chopped[2][7] = 16'b00000_110000_11111;
        rice_chopped[2][8] = 16'b00000_110000_11111;
        rice_chopped[2][9] = 16'b00000_000000_00000;
        rice_chopped[2][10] = 16'b00000_000000_00000;
        rice_chopped[2][11] = 16'b00000_000000_00000;
        rice_chopped[2][12] = 16'b00000_000000_00000;
        rice_chopped[2][13] = 16'b00000_000000_00000;
        rice_chopped[2][14] = 16'b00000_111111_00001;
        rice_chopped[3][0] = 16'b00000_111111_00001;
        rice_chopped[3][1] = 16'b00000_000000_00000;
        rice_chopped[3][2] = 16'b00000_000000_00000;
        rice_chopped[3][3] = 16'b00000_110000_11111;
        rice_chopped[3][4] = 16'b00000_110000_11111;
        rice_chopped[3][5] = 16'b00000_110000_11111;
        rice_chopped[3][6] = 16'b00000_110000_11111;
        rice_chopped[3][7] = 16'b00000_110000_11111;
        rice_chopped[3][8] = 16'b00000_110000_11111;
        rice_chopped[3][9] = 16'b00000_110000_11111;
        rice_chopped[3][10] = 16'b00000_110000_11111;
        rice_chopped[3][11] = 16'b00000_110000_11111;
        rice_chopped[3][12] = 16'b00000_000000_00000;
        rice_chopped[3][13] = 16'b00000_000000_00000;
        rice_chopped[3][14] = 16'b00000_111111_00001;
        rice_chopped[4][0] = 16'b00000_111111_00001;
        rice_chopped[4][1] = 16'b00000_000000_00000;
        rice_chopped[4][2] = 16'b00000_000000_00000;
        rice_chopped[4][3] = 16'b00000_110000_11111;
        rice_chopped[4][4] = 16'b00000_110000_11111;
        rice_chopped[4][5] = 16'b00000_110000_11111;
        rice_chopped[4][6] = 16'b00000_110000_11111;
        rice_chopped[4][7] = 16'b00000_110000_11111;
        rice_chopped[4][8] = 16'b00000_110000_11111;
        rice_chopped[4][9] = 16'b00000_110000_11111;
        rice_chopped[4][10] = 16'b00000_110000_11111;
        rice_chopped[4][11] = 16'b00000_110000_11111;
        rice_chopped[4][12] = 16'b00000_000000_00000;
        rice_chopped[4][13] = 16'b00000_000000_00000;
        rice_chopped[4][14] = 16'b00000_111111_00001;
        rice_chopped[5][0] = 16'b00000_111111_00001;
        rice_chopped[5][1] = 16'b00000_000000_00000;
        rice_chopped[5][2] = 16'b00000_110000_11111;
        rice_chopped[5][3] = 16'b00000_110000_11111;
        rice_chopped[5][4] = 16'b00000_110000_11111;
        rice_chopped[5][5] = 16'b00000_110000_11111;
        rice_chopped[5][6] = 16'b00000_110000_11111;
        rice_chopped[5][7] = 16'b00000_110000_11111;
        rice_chopped[5][8] = 16'b00000_110000_11111;
        rice_chopped[5][9] = 16'b00000_110000_11111;
        rice_chopped[5][10] = 16'b00000_110000_11111;
        rice_chopped[5][11] = 16'b00000_110000_11111;
        rice_chopped[5][12] = 16'b00000_110000_11111;
        rice_chopped[5][13] = 16'b00000_000000_00000;
        rice_chopped[5][14] = 16'b00000_111111_00001;
        rice_chopped[6][0] = 16'b00000_111111_00001;
        rice_chopped[6][1] = 16'b00000_000000_00000;
        rice_chopped[6][2] = 16'b00000_110000_11111;
        rice_chopped[6][3] = 16'b00000_110000_11111;
        rice_chopped[6][4] = 16'b11111_111110_11111;
        rice_chopped[6][5] = 16'b11111_111110_11111;
        rice_chopped[6][6] = 16'b10001_100011_10001;
        rice_chopped[6][7] = 16'b11111_111110_11111;
        rice_chopped[6][8] = 16'b11111_111110_11111;
        rice_chopped[6][9] = 16'b11111_111110_11111;
        rice_chopped[6][10] = 16'b11111_111110_11111;
        rice_chopped[6][11] = 16'b00000_110000_11111;
        rice_chopped[6][12] = 16'b00000_110000_11111;
        rice_chopped[6][13] = 16'b00000_000000_00000;
        rice_chopped[6][14] = 16'b00000_111111_00001;
        rice_chopped[7][0] = 16'b00000_111111_00001;
        rice_chopped[7][1] = 16'b00000_000000_00000;
        rice_chopped[7][2] = 16'b00000_110000_11111;
        rice_chopped[7][3] = 16'b11111_111110_11111;
        rice_chopped[7][4] = 16'b11111_111110_11111;
        rice_chopped[7][5] = 16'b11111_111110_11111;
        rice_chopped[7][6] = 16'b11111_111110_11111;
        rice_chopped[7][7] = 16'b11111_111110_11111;
        rice_chopped[7][8] = 16'b11111_111110_11111;
        rice_chopped[7][9] = 16'b10001_100011_10001;
        rice_chopped[7][10] = 16'b11111_111110_11111;
        rice_chopped[7][11] = 16'b11111_111110_11111;
        rice_chopped[7][12] = 16'b00000_110000_11111;
        rice_chopped[7][13] = 16'b00000_000000_00000;
        rice_chopped[7][14] = 16'b00000_111111_00001;
        rice_chopped[8][0] = 16'b00000_111111_00001;
        rice_chopped[8][1] = 16'b00000_000000_00000;
        rice_chopped[8][2] = 16'b00000_000000_00000;
        rice_chopped[8][3] = 16'b10001_100011_10001;
        rice_chopped[8][4] = 16'b11111_111110_11111;
        rice_chopped[8][5] = 16'b10001_100011_10001;
        rice_chopped[8][6] = 16'b11111_111110_11111;
        rice_chopped[8][7] = 16'b10001_100011_10001;
        rice_chopped[8][8] = 16'b11111_111110_11111;
        rice_chopped[8][9] = 16'b11111_111110_11111;
        rice_chopped[8][10] = 16'b11111_111110_11111;
        rice_chopped[8][11] = 16'b10001_100011_10001;
        rice_chopped[8][12] = 16'b00000_000000_00000;
        rice_chopped[8][13] = 16'b00000_000000_00000;
        rice_chopped[8][14] = 16'b00000_111111_00001;
        rice_chopped[9][0] = 16'b00000_111111_00001;
        rice_chopped[9][1] = 16'b00000_000000_00000;
        rice_chopped[9][2] = 16'b00000_000000_00000;
        rice_chopped[9][3] = 16'b11111_111110_11111;
        rice_chopped[9][4] = 16'b11111_111110_11111;
        rice_chopped[9][5] = 16'b11111_111110_11111;
        rice_chopped[9][6] = 16'b11111_111110_11111;
        rice_chopped[9][7] = 16'b11111_111110_11111;
        rice_chopped[9][8] = 16'b11111_111110_11111;
        rice_chopped[9][9] = 16'b10001_100011_10001;
        rice_chopped[9][10] = 16'b11111_111110_11111;
        rice_chopped[9][11] = 16'b11111_111110_11111;
        rice_chopped[9][12] = 16'b00000_000000_00000;
        rice_chopped[9][13] = 16'b00000_000000_00000;
        rice_chopped[9][14] = 16'b00000_111111_00001;
        rice_chopped[10][0] = 16'b00000_111111_00001;
        rice_chopped[10][1] = 16'b00000_000000_00000;
        rice_chopped[10][2] = 16'b00000_000000_00000;
        rice_chopped[10][3] = 16'b00000_000000_00000;
        rice_chopped[10][4] = 16'b11111_111110_11111;
        rice_chopped[10][5] = 16'b11111_111110_11111;
        rice_chopped[10][6] = 16'b10001_100011_10001;
        rice_chopped[10][7] = 16'b11111_111110_11111;
        rice_chopped[10][8] = 16'b11111_111110_11111;
        rice_chopped[10][9] = 16'b11111_111110_11111;
        rice_chopped[10][10] = 16'b11111_111110_11111;
        rice_chopped[10][11] = 16'b00000_000000_00000;
        rice_chopped[10][12] = 16'b00000_000000_00000;
        rice_chopped[10][13] = 16'b00000_000000_00000;
        rice_chopped[10][14] = 16'b00000_111111_00001;
        rice_chopped[11][0] = 16'b00000_111111_00001;
        rice_chopped[11][1] = 16'b00000_000000_00000;
        rice_chopped[11][2] = 16'b00000_000000_00000;
        rice_chopped[11][3] = 16'b00000_000000_00000;
        rice_chopped[11][4] = 16'b00000_000000_00000;
        rice_chopped[11][5] = 16'b11111_111110_11111;
        rice_chopped[11][6] = 16'b11111_111110_11111;
        rice_chopped[11][7] = 16'b11111_111110_11111;
        rice_chopped[11][8] = 16'b10001_100011_10001;
        rice_chopped[11][9] = 16'b11111_111110_11111;
        rice_chopped[11][10] = 16'b00000_000000_00000;
        rice_chopped[11][11] = 16'b00000_000000_00000;
        rice_chopped[11][12] = 16'b00000_000000_00000;
        rice_chopped[11][13] = 16'b00000_000000_00000;
        rice_chopped[11][14] = 16'b00000_111111_00001;
        rice_chopped[12][0] = 16'b00000_111111_00001;
        rice_chopped[12][1] = 16'b00000_000000_00000;
        rice_chopped[12][2] = 16'b00000_000000_00000;
        rice_chopped[12][3] = 16'b00000_000000_00000;
        rice_chopped[12][4] = 16'b00000_000000_00000;
        rice_chopped[12][5] = 16'b00000_000000_00000;
        rice_chopped[12][6] = 16'b11111_111110_11111;
        rice_chopped[12][7] = 16'b11111_111110_11111;
        rice_chopped[12][8] = 16'b11111_111110_11111;
        rice_chopped[12][9] = 16'b00000_000000_00000;
        rice_chopped[12][10] = 16'b00000_000000_00000;
        rice_chopped[12][11] = 16'b00000_000000_00000;
        rice_chopped[12][12] = 16'b00000_000000_00000;
        rice_chopped[12][13] = 16'b00000_000000_00000;
        rice_chopped[12][14] = 16'b00000_111111_00001;
        rice_chopped[13][0] = 16'b00000_111111_00001;
        rice_chopped[13][1] = 16'b00000_000000_00000;
        rice_chopped[13][2] = 16'b00000_000000_00000;
        rice_chopped[13][3] = 16'b00000_000000_00000;
        rice_chopped[13][4] = 16'b00000_000000_00000;
        rice_chopped[13][5] = 16'b00000_000000_00000;
        rice_chopped[13][6] = 16'b00000_000000_00000;
        rice_chopped[13][7] = 16'b00000_000000_00000;
        rice_chopped[13][8] = 16'b00000_000000_00000;
        rice_chopped[13][9] = 16'b00000_000000_00000;
        rice_chopped[13][10] = 16'b00000_000000_00000;
        rice_chopped[13][11] = 16'b00000_000000_00000;
        rice_chopped[13][12] = 16'b00000_000000_00000;
        rice_chopped[13][13] = 16'b00000_000000_00000;
        rice_chopped[13][14] = 16'b00000_111111_00001;
        rice_chopped[14][0] = 16'b00000_111111_00001;
        rice_chopped[14][1] = 16'b00000_111111_00001;
        rice_chopped[14][2] = 16'b00000_111111_00001;
        rice_chopped[14][3] = 16'b00000_111111_00001;
        rice_chopped[14][4] = 16'b00000_111111_00001;
        rice_chopped[14][5] = 16'b00000_111111_00001;
        rice_chopped[14][6] = 16'b00000_111111_00001;
        rice_chopped[14][7] = 16'b00000_111111_00001;
        rice_chopped[14][8] = 16'b00000_111111_00001;
        rice_chopped[14][9] = 16'b00000_111111_00001;
        rice_chopped[14][10] = 16'b00000_111111_00001;
        rice_chopped[14][11] = 16'b00000_111111_00001;
        rice_chopped[14][12] = 16'b00000_111111_00001;
        rice_chopped[14][13] = 16'b00000_111111_00001;
        rice_chopped[14][14] = 16'b00000_111111_00001;

        
        rice_boiled_chopped[0][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][1] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][2] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][3] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][4] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][5] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][6] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][7] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][8] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][9] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][10] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][11] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][12] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][13] = 16'b10101_011000_00000;
        rice_boiled_chopped[0][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[1][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[1][1] = 16'b00000_000000_00000;
        rice_boiled_chopped[1][2] = 16'b00000_000000_00000;
        rice_boiled_chopped[1][3] = 16'b00000_000000_00000;
        rice_boiled_chopped[1][4] = 16'b00000_000000_00000;
        rice_boiled_chopped[1][5] = 16'b00000_000000_00000;
        rice_boiled_chopped[1][6] = 16'b00000_000000_00000;
        rice_boiled_chopped[1][7] = 16'b00000_000000_00000;
        rice_boiled_chopped[1][8] = 16'b00000_000000_00000;
        rice_boiled_chopped[1][9] = 16'b00000_000000_00000;
        rice_boiled_chopped[1][10] = 16'b00000_000000_00000;
        rice_boiled_chopped[1][11] = 16'b00000_000000_00000;
        rice_boiled_chopped[1][12] = 16'b00000_000000_00000;
        rice_boiled_chopped[1][13] = 16'b00000_000000_00000;
        rice_boiled_chopped[1][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[2][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[2][1] = 16'b00000_000000_00000;
        rice_boiled_chopped[2][2] = 16'b00000_000000_00000;
        rice_boiled_chopped[2][3] = 16'b00000_000000_00000;
        rice_boiled_chopped[2][4] = 16'b00000_000000_00000;
        rice_boiled_chopped[2][5] = 16'b00000_000000_00000;
        rice_boiled_chopped[2][6] = 16'b00000_110000_11111;
        rice_boiled_chopped[2][7] = 16'b00000_110000_11111;
        rice_boiled_chopped[2][8] = 16'b00000_110000_11111;
        rice_boiled_chopped[2][9] = 16'b00000_000000_00000;
        rice_boiled_chopped[2][10] = 16'b00000_000000_00000;
        rice_boiled_chopped[2][11] = 16'b00000_000000_00000;
        rice_boiled_chopped[2][12] = 16'b00000_000000_00000;
        rice_boiled_chopped[2][13] = 16'b00000_000000_00000;
        rice_boiled_chopped[2][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[3][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[3][1] = 16'b00000_000000_00000;
        rice_boiled_chopped[3][2] = 16'b00000_000000_00000;
        rice_boiled_chopped[3][3] = 16'b00000_110000_11111;
        rice_boiled_chopped[3][4] = 16'b00000_110000_11111;
        rice_boiled_chopped[3][5] = 16'b00000_110000_11111;
        rice_boiled_chopped[3][6] = 16'b00000_110000_11111;
        rice_boiled_chopped[3][7] = 16'b00000_110000_11111;
        rice_boiled_chopped[3][8] = 16'b00000_110000_11111;
        rice_boiled_chopped[3][9] = 16'b00000_110000_11111;
        rice_boiled_chopped[3][10] = 16'b00000_110000_11111;
        rice_boiled_chopped[3][11] = 16'b00000_110000_11111;
        rice_boiled_chopped[3][12] = 16'b00000_000000_00000;
        rice_boiled_chopped[3][13] = 16'b00000_000000_00000;
        rice_boiled_chopped[3][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[4][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[4][1] = 16'b00000_000000_00000;
        rice_boiled_chopped[4][2] = 16'b00000_000000_00000;
        rice_boiled_chopped[4][3] = 16'b00000_110000_11111;
        rice_boiled_chopped[4][4] = 16'b00000_110000_11111;
        rice_boiled_chopped[4][5] = 16'b00000_110000_11111;
        rice_boiled_chopped[4][6] = 16'b00000_110000_11111;
        rice_boiled_chopped[4][7] = 16'b00000_110000_11111;
        rice_boiled_chopped[4][8] = 16'b00000_110000_11111;
        rice_boiled_chopped[4][9] = 16'b00000_110000_11111;
        rice_boiled_chopped[4][10] = 16'b00000_110000_11111;
        rice_boiled_chopped[4][11] = 16'b00000_110000_11111;
        rice_boiled_chopped[4][12] = 16'b00000_000000_00000;
        rice_boiled_chopped[4][13] = 16'b00000_000000_00000;
        rice_boiled_chopped[4][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[5][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[5][1] = 16'b00000_000000_00000;
        rice_boiled_chopped[5][2] = 16'b00000_110000_11111;
        rice_boiled_chopped[5][3] = 16'b00000_110000_11111;
        rice_boiled_chopped[5][4] = 16'b00000_110000_11111;
        rice_boiled_chopped[5][5] = 16'b00000_110000_11111;
        rice_boiled_chopped[5][6] = 16'b00000_110000_11111;
        rice_boiled_chopped[5][7] = 16'b00000_110000_11111;
        rice_boiled_chopped[5][8] = 16'b00000_110000_11111;
        rice_boiled_chopped[5][9] = 16'b00000_110000_11111;
        rice_boiled_chopped[5][10] = 16'b00000_110000_11111;
        rice_boiled_chopped[5][11] = 16'b00000_110000_11111;
        rice_boiled_chopped[5][12] = 16'b00000_110000_11111;
        rice_boiled_chopped[5][13] = 16'b00000_000000_00000;
        rice_boiled_chopped[5][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[6][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[6][1] = 16'b00000_000000_00000;
        rice_boiled_chopped[6][2] = 16'b00000_110000_11111;
        rice_boiled_chopped[6][3] = 16'b00000_110000_11111;
        rice_boiled_chopped[6][4] = 16'b11111_111110_11111;
        rice_boiled_chopped[6][5] = 16'b11111_111110_11111;
        rice_boiled_chopped[6][6] = 16'b10001_100011_10001;
        rice_boiled_chopped[6][7] = 16'b11111_111110_11111;
        rice_boiled_chopped[6][8] = 16'b11111_111110_11111;
        rice_boiled_chopped[6][9] = 16'b11111_111110_11111;
        rice_boiled_chopped[6][10] = 16'b11111_111110_11111;
        rice_boiled_chopped[6][11] = 16'b00000_110000_11111;
        rice_boiled_chopped[6][12] = 16'b00000_110000_11111;
        rice_boiled_chopped[6][13] = 16'b00000_000000_00000;
        rice_boiled_chopped[6][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[7][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[7][1] = 16'b00000_000000_00000;
        rice_boiled_chopped[7][2] = 16'b00000_110000_11111;
        rice_boiled_chopped[7][3] = 16'b11111_111110_11111;
        rice_boiled_chopped[7][4] = 16'b11111_111110_11111;
        rice_boiled_chopped[7][5] = 16'b11111_111110_11111;
        rice_boiled_chopped[7][6] = 16'b11111_111110_11111;
        rice_boiled_chopped[7][7] = 16'b11111_111110_11111;
        rice_boiled_chopped[7][8] = 16'b11111_111110_11111;
        rice_boiled_chopped[7][9] = 16'b10001_100011_10001;
        rice_boiled_chopped[7][10] = 16'b11111_111110_11111;
        rice_boiled_chopped[7][11] = 16'b11111_111110_11111;
        rice_boiled_chopped[7][12] = 16'b00000_110000_11111;
        rice_boiled_chopped[7][13] = 16'b00000_000000_00000;
        rice_boiled_chopped[7][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[8][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[8][1] = 16'b00000_000000_00000;
        rice_boiled_chopped[8][2] = 16'b00000_000000_00000;
        rice_boiled_chopped[8][3] = 16'b10001_100011_10001;
        rice_boiled_chopped[8][4] = 16'b11111_111110_11111;
        rice_boiled_chopped[8][5] = 16'b10001_100011_10001;
        rice_boiled_chopped[8][6] = 16'b11111_111110_11111;
        rice_boiled_chopped[8][7] = 16'b10001_100011_10001;
        rice_boiled_chopped[8][8] = 16'b11111_111110_11111;
        rice_boiled_chopped[8][9] = 16'b11111_111110_11111;
        rice_boiled_chopped[8][10] = 16'b11111_111110_11111;
        rice_boiled_chopped[8][11] = 16'b10001_100011_10001;
        rice_boiled_chopped[8][12] = 16'b00000_000000_00000;
        rice_boiled_chopped[8][13] = 16'b00000_000000_00000;
        rice_boiled_chopped[8][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[9][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[9][1] = 16'b00000_000000_00000;
        rice_boiled_chopped[9][2] = 16'b00000_000000_00000;
        rice_boiled_chopped[9][3] = 16'b11111_111110_11111;
        rice_boiled_chopped[9][4] = 16'b11111_111110_11111;
        rice_boiled_chopped[9][5] = 16'b11111_111110_11111;
        rice_boiled_chopped[9][6] = 16'b11111_111110_11111;
        rice_boiled_chopped[9][7] = 16'b11111_111110_11111;
        rice_boiled_chopped[9][8] = 16'b11111_111110_11111;
        rice_boiled_chopped[9][9] = 16'b10001_100011_10001;
        rice_boiled_chopped[9][10] = 16'b11111_111110_11111;
        rice_boiled_chopped[9][11] = 16'b11111_111110_11111;
        rice_boiled_chopped[9][12] = 16'b00000_000000_00000;
        rice_boiled_chopped[9][13] = 16'b00000_000000_00000;
        rice_boiled_chopped[9][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[10][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[10][1] = 16'b00000_000000_00000;
        rice_boiled_chopped[10][2] = 16'b00000_000000_00000;
        rice_boiled_chopped[10][3] = 16'b00000_000000_00000;
        rice_boiled_chopped[10][4] = 16'b11111_111110_11111;
        rice_boiled_chopped[10][5] = 16'b11111_111110_11111;
        rice_boiled_chopped[10][6] = 16'b10001_100011_10001;
        rice_boiled_chopped[10][7] = 16'b11111_111110_11111;
        rice_boiled_chopped[10][8] = 16'b11111_111110_11111;
        rice_boiled_chopped[10][9] = 16'b11111_111110_11111;
        rice_boiled_chopped[10][10] = 16'b11111_111110_11111;
        rice_boiled_chopped[10][11] = 16'b00000_000000_00000;
        rice_boiled_chopped[10][12] = 16'b00000_000000_00000;
        rice_boiled_chopped[10][13] = 16'b00000_000000_00000;
        rice_boiled_chopped[10][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[11][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[11][1] = 16'b00000_000000_00000;
        rice_boiled_chopped[11][2] = 16'b00000_000000_00000;
        rice_boiled_chopped[11][3] = 16'b00000_000000_00000;
        rice_boiled_chopped[11][4] = 16'b00000_000000_00000;
        rice_boiled_chopped[11][5] = 16'b11111_111110_11111;
        rice_boiled_chopped[11][6] = 16'b11111_111110_11111;
        rice_boiled_chopped[11][7] = 16'b11111_111110_11111;
        rice_boiled_chopped[11][8] = 16'b10001_100011_10001;
        rice_boiled_chopped[11][9] = 16'b11111_111110_11111;
        rice_boiled_chopped[11][10] = 16'b00000_000000_00000;
        rice_boiled_chopped[11][11] = 16'b00000_000000_00000;
        rice_boiled_chopped[11][12] = 16'b00000_000000_00000;
        rice_boiled_chopped[11][13] = 16'b00000_000000_00000;
        rice_boiled_chopped[11][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[12][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[12][1] = 16'b00000_000000_00000;
        rice_boiled_chopped[12][2] = 16'b00000_000000_00000;
        rice_boiled_chopped[12][3] = 16'b00000_000000_00000;
        rice_boiled_chopped[12][4] = 16'b00000_000000_00000;
        rice_boiled_chopped[12][5] = 16'b00000_000000_00000;
        rice_boiled_chopped[12][6] = 16'b11111_111110_11111;
        rice_boiled_chopped[12][7] = 16'b11111_111110_11111;
        rice_boiled_chopped[12][8] = 16'b11111_111110_11111;
        rice_boiled_chopped[12][9] = 16'b00000_000000_00000;
        rice_boiled_chopped[12][10] = 16'b00000_000000_00000;
        rice_boiled_chopped[12][11] = 16'b00000_000000_00000;
        rice_boiled_chopped[12][12] = 16'b00000_000000_00000;
        rice_boiled_chopped[12][13] = 16'b00000_000000_00000;
        rice_boiled_chopped[12][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[13][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[13][1] = 16'b00000_000000_00000;
        rice_boiled_chopped[13][2] = 16'b00000_000000_00000;
        rice_boiled_chopped[13][3] = 16'b00000_000000_00000;
        rice_boiled_chopped[13][4] = 16'b00000_000000_00000;
        rice_boiled_chopped[13][5] = 16'b00000_000000_00000;
        rice_boiled_chopped[13][6] = 16'b00000_000000_00000;
        rice_boiled_chopped[13][7] = 16'b00000_000000_00000;
        rice_boiled_chopped[13][8] = 16'b00000_000000_00000;
        rice_boiled_chopped[13][9] = 16'b00000_000000_00000;
        rice_boiled_chopped[13][10] = 16'b00000_000000_00000;
        rice_boiled_chopped[13][11] = 16'b00000_000000_00000;
        rice_boiled_chopped[13][12] = 16'b00000_000000_00000;
        rice_boiled_chopped[13][13] = 16'b00000_000000_00000;
        rice_boiled_chopped[13][14] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][0] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][1] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][2] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][3] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][4] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][5] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][6] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][7] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][8] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][9] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][10] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][11] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][12] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][13] = 16'b10101_011000_00000;
        rice_boiled_chopped[14][14] = 16'b10101_011000_00000;

        chicken_boiled_chopped[0][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][1] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][2] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][3] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][4] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][5] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][6] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][7] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][8] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][9] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][10] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][11] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][12] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][13] = 16'b10101_011000_00000;
        chicken_boiled_chopped[0][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[1][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[1][1] = 16'b11111_111110_11111;
        chicken_boiled_chopped[1][2] = 16'b11111_111110_11111;
        chicken_boiled_chopped[1][3] = 16'b00000_000000_00000;
        chicken_boiled_chopped[1][4] = 16'b00000_000000_00000;
        chicken_boiled_chopped[1][5] = 16'b00000_000000_00000;
        chicken_boiled_chopped[1][6] = 16'b00000_000000_00000;
        chicken_boiled_chopped[1][7] = 16'b00000_000000_00000;
        chicken_boiled_chopped[1][8] = 16'b00000_000000_00000;
        chicken_boiled_chopped[1][9] = 16'b00000_000000_00000;
        chicken_boiled_chopped[1][10] = 16'b00000_000000_00000;
        chicken_boiled_chopped[1][11] = 16'b00000_000000_00000;
        chicken_boiled_chopped[1][12] = 16'b00000_000000_00000;
        chicken_boiled_chopped[1][13] = 16'b00000_000000_00000;
        chicken_boiled_chopped[1][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[2][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[2][1] = 16'b11111_111110_11111;
        chicken_boiled_chopped[2][2] = 16'b11111_111110_11111;
        chicken_boiled_chopped[2][3] = 16'b11111_111110_11111;
        chicken_boiled_chopped[2][4] = 16'b00000_000000_00000;
        chicken_boiled_chopped[2][5] = 16'b00000_000000_00000;
        chicken_boiled_chopped[2][6] = 16'b00000_000000_00000;
        chicken_boiled_chopped[2][7] = 16'b00000_000000_00000;
        chicken_boiled_chopped[2][8] = 16'b00000_000000_00000;
        chicken_boiled_chopped[2][9] = 16'b00000_000000_00000;
        chicken_boiled_chopped[2][10] = 16'b00000_000000_00000;
        chicken_boiled_chopped[2][11] = 16'b00000_000000_00000;
        chicken_boiled_chopped[2][12] = 16'b00000_000000_00000;
        chicken_boiled_chopped[2][13] = 16'b00000_000000_00000;
        chicken_boiled_chopped[2][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[3][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[3][1] = 16'b00000_000000_00000;
        chicken_boiled_chopped[3][2] = 16'b11111_111110_11111;
        chicken_boiled_chopped[3][3] = 16'b11111_111110_11111;
        chicken_boiled_chopped[3][4] = 16'b11111_111110_11111;
        chicken_boiled_chopped[3][5] = 16'b00000_000000_00000;
        chicken_boiled_chopped[3][6] = 16'b00000_000000_00000;
        chicken_boiled_chopped[3][7] = 16'b00000_000000_00000;
        chicken_boiled_chopped[3][8] = 16'b00000_000000_00000;
        chicken_boiled_chopped[3][9] = 16'b00000_000000_00000;
        chicken_boiled_chopped[3][10] = 16'b00000_000000_00000;
        chicken_boiled_chopped[3][11] = 16'b00000_000000_00000;
        chicken_boiled_chopped[3][12] = 16'b00000_000000_00000;
        chicken_boiled_chopped[3][13] = 16'b00000_000000_00000;
        chicken_boiled_chopped[3][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[4][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[4][1] = 16'b00000_000000_00000;
        chicken_boiled_chopped[4][2] = 16'b00000_000000_00000;
        chicken_boiled_chopped[4][3] = 16'b11111_111110_11111;
        chicken_boiled_chopped[4][4] = 16'b11111_101000_00100;
        chicken_boiled_chopped[4][5] = 16'b11111_101000_00100;
        chicken_boiled_chopped[4][6] = 16'b11111_101000_00100;
        chicken_boiled_chopped[4][7] = 16'b00000_000000_00000;
        chicken_boiled_chopped[4][8] = 16'b00000_000000_00000;
        chicken_boiled_chopped[4][9] = 16'b00000_000000_00000;
        chicken_boiled_chopped[4][10] = 16'b00000_000000_00000;
        chicken_boiled_chopped[4][11] = 16'b00000_000000_00000;
        chicken_boiled_chopped[4][12] = 16'b00000_000000_00000;
        chicken_boiled_chopped[4][13] = 16'b00000_000000_00000;
        chicken_boiled_chopped[4][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[5][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[5][1] = 16'b00000_000000_00000;
        chicken_boiled_chopped[5][2] = 16'b00000_000000_00000;
        chicken_boiled_chopped[5][3] = 16'b00000_000000_00000;
        chicken_boiled_chopped[5][4] = 16'b11111_101000_00100;
        chicken_boiled_chopped[5][5] = 16'b11111_101111_01111;
        chicken_boiled_chopped[5][6] = 16'b11111_101111_01111;
        chicken_boiled_chopped[5][7] = 16'b11111_101000_00100;
        chicken_boiled_chopped[5][8] = 16'b11111_101000_00100;
        chicken_boiled_chopped[5][9] = 16'b00000_000000_00000;
        chicken_boiled_chopped[5][10] = 16'b00000_000000_00000;
        chicken_boiled_chopped[5][11] = 16'b00000_000000_00000;
        chicken_boiled_chopped[5][12] = 16'b00000_000000_00000;
        chicken_boiled_chopped[5][13] = 16'b00000_000000_00000;
        chicken_boiled_chopped[5][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[6][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[6][1] = 16'b00000_000000_00000;
        chicken_boiled_chopped[6][2] = 16'b00000_000000_00000;
        chicken_boiled_chopped[6][3] = 16'b00000_000000_00000;
        chicken_boiled_chopped[6][4] = 16'b00000_000000_00000;
        chicken_boiled_chopped[6][5] = 16'b11111_101000_00100;
        chicken_boiled_chopped[6][6] = 16'b11111_101111_01111;
        chicken_boiled_chopped[6][7] = 16'b11111_101111_01111;
        chicken_boiled_chopped[6][8] = 16'b11111_101111_01111;
        chicken_boiled_chopped[6][9] = 16'b11111_101000_00100;
        chicken_boiled_chopped[6][10] = 16'b11111_101000_00100;
        chicken_boiled_chopped[6][11] = 16'b11111_101000_00100;
        chicken_boiled_chopped[6][12] = 16'b00000_000000_00000;
        chicken_boiled_chopped[6][13] = 16'b00000_000000_00000;
        chicken_boiled_chopped[6][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[7][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[7][1] = 16'b00000_000000_00000;
        chicken_boiled_chopped[7][2] = 16'b00000_000000_00000;
        chicken_boiled_chopped[7][3] = 16'b00000_000000_00000;
        chicken_boiled_chopped[7][4] = 16'b00000_000000_00000;
        chicken_boiled_chopped[7][5] = 16'b11111_101000_00100;
        chicken_boiled_chopped[7][6] = 16'b11111_101111_01111;
        chicken_boiled_chopped[7][7] = 16'b11111_101111_01111;
        chicken_boiled_chopped[7][8] = 16'b11111_101111_01111;
        chicken_boiled_chopped[7][9] = 16'b11111_101111_01111;
        chicken_boiled_chopped[7][10] = 16'b11111_101111_01111;
        chicken_boiled_chopped[7][11] = 16'b11111_101000_00100;
        chicken_boiled_chopped[7][12] = 16'b11111_101000_00100;
        chicken_boiled_chopped[7][13] = 16'b00000_000000_00000;
        chicken_boiled_chopped[7][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[8][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[8][1] = 16'b00000_000000_00000;
        chicken_boiled_chopped[8][2] = 16'b00000_000000_00000;
        chicken_boiled_chopped[8][3] = 16'b00000_000000_00000;
        chicken_boiled_chopped[8][4] = 16'b00000_000000_00000;
        chicken_boiled_chopped[8][5] = 16'b00000_000000_00000;
        chicken_boiled_chopped[8][6] = 16'b11111_101000_00100;
        chicken_boiled_chopped[8][7] = 16'b11111_101111_01111;
        chicken_boiled_chopped[8][8] = 16'b11111_101111_01111;
        chicken_boiled_chopped[8][9] = 16'b11111_101111_01111;
        chicken_boiled_chopped[8][10] = 16'b11111_101111_01111;
        chicken_boiled_chopped[8][11] = 16'b11111_101111_01111;
        chicken_boiled_chopped[8][12] = 16'b11111_101000_00100;
        chicken_boiled_chopped[8][13] = 16'b00000_000000_00000;
        chicken_boiled_chopped[8][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[9][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[9][1] = 16'b00000_000000_00000;
        chicken_boiled_chopped[9][2] = 16'b00000_000000_00000;
        chicken_boiled_chopped[9][3] = 16'b00000_000000_00000;
        chicken_boiled_chopped[9][4] = 16'b00000_000000_00000;
        chicken_boiled_chopped[9][5] = 16'b00000_000000_00000;
        chicken_boiled_chopped[9][6] = 16'b11111_101000_00100;
        chicken_boiled_chopped[9][7] = 16'b11111_101111_01111;
        chicken_boiled_chopped[9][8] = 16'b11111_101111_01111;
        chicken_boiled_chopped[9][9] = 16'b11111_101111_01111;
        chicken_boiled_chopped[9][10] = 16'b11111_101111_01111;
        chicken_boiled_chopped[9][11] = 16'b11111_101111_01111;
        chicken_boiled_chopped[9][12] = 16'b11111_101000_00100;
        chicken_boiled_chopped[9][13] = 16'b11111_101000_00100;
        chicken_boiled_chopped[9][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[10][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[10][1] = 16'b00000_000000_00000;
        chicken_boiled_chopped[10][2] = 16'b00000_000000_00000;
        chicken_boiled_chopped[10][3] = 16'b00000_000000_00000;
        chicken_boiled_chopped[10][4] = 16'b00000_000000_00000;
        chicken_boiled_chopped[10][5] = 16'b00000_000000_00000;
        chicken_boiled_chopped[10][6] = 16'b11111_101000_00100;
        chicken_boiled_chopped[10][7] = 16'b11111_101111_01111;
        chicken_boiled_chopped[10][8] = 16'b11111_101111_01111;
        chicken_boiled_chopped[10][9] = 16'b11111_101111_01111;
        chicken_boiled_chopped[10][10] = 16'b11111_101111_01111;
        chicken_boiled_chopped[10][11] = 16'b11111_101111_01111;
        chicken_boiled_chopped[10][12] = 16'b11111_101111_01111;
        chicken_boiled_chopped[10][13] = 16'b11111_101000_00100;
        chicken_boiled_chopped[10][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[11][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[11][1] = 16'b00000_000000_00000;
        chicken_boiled_chopped[11][2] = 16'b00000_000000_00000;
        chicken_boiled_chopped[11][3] = 16'b00000_000000_00000;
        chicken_boiled_chopped[11][4] = 16'b00000_000000_00000;
        chicken_boiled_chopped[11][5] = 16'b00000_000000_00000;
        chicken_boiled_chopped[11][6] = 16'b00000_000000_00000;
        chicken_boiled_chopped[11][7] = 16'b11111_101000_00100;
        chicken_boiled_chopped[11][8] = 16'b11111_101111_01111;
        chicken_boiled_chopped[11][9] = 16'b11111_101111_01111;
        chicken_boiled_chopped[11][10] = 16'b11111_101111_01111;
        chicken_boiled_chopped[11][11] = 16'b11111_101111_01111;
        chicken_boiled_chopped[11][12] = 16'b11111_101000_00100;
        chicken_boiled_chopped[11][13] = 16'b11111_101000_00100;
        chicken_boiled_chopped[11][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[12][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[12][1] = 16'b00000_000000_00000;
        chicken_boiled_chopped[12][2] = 16'b00000_000000_00000;
        chicken_boiled_chopped[12][3] = 16'b00000_000000_00000;
        chicken_boiled_chopped[12][4] = 16'b00000_000000_00000;
        chicken_boiled_chopped[12][5] = 16'b00000_000000_00000;
        chicken_boiled_chopped[12][6] = 16'b00000_000000_00000;
        chicken_boiled_chopped[12][7] = 16'b11111_101000_00100;
        chicken_boiled_chopped[12][8] = 16'b11111_101000_00100;
        chicken_boiled_chopped[12][9] = 16'b11111_101111_01111;
        chicken_boiled_chopped[12][10] = 16'b11111_101111_01111;
        chicken_boiled_chopped[12][11] = 16'b11111_101111_01111;
        chicken_boiled_chopped[12][12] = 16'b11111_101000_00100;
        chicken_boiled_chopped[12][13] = 16'b00000_000000_00000;
        chicken_boiled_chopped[12][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[13][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[13][1] = 16'b00000_000000_00000;
        chicken_boiled_chopped[13][2] = 16'b00000_000000_00000;
        chicken_boiled_chopped[13][3] = 16'b00000_000000_00000;
        chicken_boiled_chopped[13][4] = 16'b00000_000000_00000;
        chicken_boiled_chopped[13][5] = 16'b00000_000000_00000;
        chicken_boiled_chopped[13][6] = 16'b00000_000000_00000;
        chicken_boiled_chopped[13][7] = 16'b00000_000000_00000;
        chicken_boiled_chopped[13][8] = 16'b00000_000000_00000;
        chicken_boiled_chopped[13][9] = 16'b11111_101000_00100;
        chicken_boiled_chopped[13][10] = 16'b11111_101000_00100;
        chicken_boiled_chopped[13][11] = 16'b11111_101000_00100;
        chicken_boiled_chopped[13][12] = 16'b00000_000000_00000;
        chicken_boiled_chopped[13][13] = 16'b00000_000000_00000;
        chicken_boiled_chopped[13][14] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][0] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][1] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][2] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][3] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][4] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][5] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][6] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][7] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][8] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][9] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][10] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][11] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][12] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][13] = 16'b10101_011000_00000;
        chicken_boiled_chopped[14][14] = 16'b10101_011000_00000;


        chicken_boiled[0][0] = 16'b00000_000110_11111;
        chicken_boiled[0][1] = 16'b00000_000110_11111;
        chicken_boiled[0][2] = 16'b00000_000110_11111;
        chicken_boiled[0][3] = 16'b00000_000110_11111;
        chicken_boiled[0][4] = 16'b00000_000110_11111;
        chicken_boiled[0][5] = 16'b00000_000110_11111;
        chicken_boiled[0][6] = 16'b00000_000110_11111;
        chicken_boiled[0][7] = 16'b00000_000110_11111;
        chicken_boiled[0][8] = 16'b00000_000110_11111;
        chicken_boiled[0][9] = 16'b00000_000110_11111;
        chicken_boiled[0][10] = 16'b00000_000110_11111;
        chicken_boiled[0][11] = 16'b00000_000110_11111;
        chicken_boiled[0][12] = 16'b00000_000110_11111;
        chicken_boiled[0][13] = 16'b00000_000110_11111;
        chicken_boiled[0][14] = 16'b00000_000110_11111;
        chicken_boiled[1][0] = 16'b00000_000110_11111;
        chicken_boiled[1][1] = 16'b11111_111110_11111;
        chicken_boiled[1][2] = 16'b11111_111110_11111;
        chicken_boiled[1][3] = 16'b00000_000000_00000;
        chicken_boiled[1][4] = 16'b00000_000000_00000;
        chicken_boiled[1][5] = 16'b00000_000000_00000;
        chicken_boiled[1][6] = 16'b00000_000000_00000;
        chicken_boiled[1][7] = 16'b00000_000000_00000;
        chicken_boiled[1][8] = 16'b00000_000000_00000;
        chicken_boiled[1][9] = 16'b00000_000000_00000;
        chicken_boiled[1][10] = 16'b00000_000000_00000;
        chicken_boiled[1][11] = 16'b00000_000000_00000;
        chicken_boiled[1][12] = 16'b00000_000000_00000;
        chicken_boiled[1][13] = 16'b00000_000000_00000;
        chicken_boiled[1][14] = 16'b00000_000110_11111;
        chicken_boiled[2][0] = 16'b00000_000110_11111;
        chicken_boiled[2][1] = 16'b11111_111110_11111;
        chicken_boiled[2][2] = 16'b11111_111110_11111;
        chicken_boiled[2][3] = 16'b11111_111110_11111;
        chicken_boiled[2][4] = 16'b00000_000000_00000;
        chicken_boiled[2][5] = 16'b00000_000000_00000;
        chicken_boiled[2][6] = 16'b00000_000000_00000;
        chicken_boiled[2][7] = 16'b00000_000000_00000;
        chicken_boiled[2][8] = 16'b00000_000000_00000;
        chicken_boiled[2][9] = 16'b00000_000000_00000;
        chicken_boiled[2][10] = 16'b00000_000000_00000;
        chicken_boiled[2][11] = 16'b00000_000000_00000;
        chicken_boiled[2][12] = 16'b00000_000000_00000;
        chicken_boiled[2][13] = 16'b00000_000000_00000;
        chicken_boiled[2][14] = 16'b00000_000110_11111;
        chicken_boiled[3][0] = 16'b00000_000110_11111;
        chicken_boiled[3][1] = 16'b00000_000000_00000;
        chicken_boiled[3][2] = 16'b11111_111110_11111;
        chicken_boiled[3][3] = 16'b11111_111110_11111;
        chicken_boiled[3][4] = 16'b11111_111110_11111;
        chicken_boiled[3][5] = 16'b00000_000000_00000;
        chicken_boiled[3][6] = 16'b00000_000000_00000;
        chicken_boiled[3][7] = 16'b00000_000000_00000;
        chicken_boiled[3][8] = 16'b00000_000000_00000;
        chicken_boiled[3][9] = 16'b00000_000000_00000;
        chicken_boiled[3][10] = 16'b00000_000000_00000;
        chicken_boiled[3][11] = 16'b00000_000000_00000;
        chicken_boiled[3][12] = 16'b00000_000000_00000;
        chicken_boiled[3][13] = 16'b00000_000000_00000;
        chicken_boiled[3][14] = 16'b00000_000110_11111;
        chicken_boiled[4][0] = 16'b00000_000110_11111;
        chicken_boiled[4][1] = 16'b00000_000000_00000;
        chicken_boiled[4][2] = 16'b00000_000000_00000;
        chicken_boiled[4][3] = 16'b11111_111110_11111;
        chicken_boiled[4][4] = 16'b11111_101000_00100;
        chicken_boiled[4][5] = 16'b11111_101000_00100;
        chicken_boiled[4][6] = 16'b11111_101000_00100;
        chicken_boiled[4][7] = 16'b00000_000000_00000;
        chicken_boiled[4][8] = 16'b00000_000000_00000;
        chicken_boiled[4][9] = 16'b00000_000000_00000;
        chicken_boiled[4][10] = 16'b00000_000000_00000;
        chicken_boiled[4][11] = 16'b00000_000000_00000;
        chicken_boiled[4][12] = 16'b00000_000000_00000;
        chicken_boiled[4][13] = 16'b00000_000000_00000;
        chicken_boiled[4][14] = 16'b00000_000110_11111;
        chicken_boiled[5][0] = 16'b00000_000110_11111;
        chicken_boiled[5][1] = 16'b00000_000000_00000;
        chicken_boiled[5][2] = 16'b00000_000000_00000;
        chicken_boiled[5][3] = 16'b00000_000000_00000;
        chicken_boiled[5][4] = 16'b11111_101000_00100;
        chicken_boiled[5][5] = 16'b11111_101111_01111;
        chicken_boiled[5][6] = 16'b11111_101111_01111;
        chicken_boiled[5][7] = 16'b11111_101000_00100;
        chicken_boiled[5][8] = 16'b11111_101000_00100;
        chicken_boiled[5][9] = 16'b00000_000000_00000;
        chicken_boiled[5][10] = 16'b00000_000000_00000;
        chicken_boiled[5][11] = 16'b00000_000000_00000;
        chicken_boiled[5][12] = 16'b00000_000000_00000;
        chicken_boiled[5][13] = 16'b00000_000000_00000;
        chicken_boiled[5][14] = 16'b00000_000110_11111;
        chicken_boiled[6][0] = 16'b00000_000110_11111;
        chicken_boiled[6][1] = 16'b00000_000000_00000;
        chicken_boiled[6][2] = 16'b00000_000000_00000;
        chicken_boiled[6][3] = 16'b00000_000000_00000;
        chicken_boiled[6][4] = 16'b00000_000000_00000;
        chicken_boiled[6][5] = 16'b11111_101000_00100;
        chicken_boiled[6][6] = 16'b11111_101111_01111;
        chicken_boiled[6][7] = 16'b11111_101111_01111;
        chicken_boiled[6][8] = 16'b11111_101111_01111;
        chicken_boiled[6][9] = 16'b11111_101000_00100;
        chicken_boiled[6][10] = 16'b11111_101000_00100;
        chicken_boiled[6][11] = 16'b11111_101000_00100;
        chicken_boiled[6][12] = 16'b00000_000000_00000;
        chicken_boiled[6][13] = 16'b00000_000000_00000;
        chicken_boiled[6][14] = 16'b00000_000110_11111;
        chicken_boiled[7][0] = 16'b00000_000110_11111;
        chicken_boiled[7][1] = 16'b00000_000000_00000;
        chicken_boiled[7][2] = 16'b00000_000000_00000;
        chicken_boiled[7][3] = 16'b00000_000000_00000;
        chicken_boiled[7][4] = 16'b00000_000000_00000;
        chicken_boiled[7][5] = 16'b11111_101000_00100;
        chicken_boiled[7][6] = 16'b11111_101111_01111;
        chicken_boiled[7][7] = 16'b11111_101111_01111;
        chicken_boiled[7][8] = 16'b11111_101111_01111;
        chicken_boiled[7][9] = 16'b11111_101111_01111;
        chicken_boiled[7][10] = 16'b11111_101111_01111;
        chicken_boiled[7][11] = 16'b11111_101000_00100;
        chicken_boiled[7][12] = 16'b11111_101000_00100;
        chicken_boiled[7][13] = 16'b00000_000000_00000;
        chicken_boiled[7][14] = 16'b00000_000110_11111;
        chicken_boiled[8][0] = 16'b00000_000110_11111;
        chicken_boiled[8][1] = 16'b00000_000000_00000;
        chicken_boiled[8][2] = 16'b00000_000000_00000;
        chicken_boiled[8][3] = 16'b00000_000000_00000;
        chicken_boiled[8][4] = 16'b00000_000000_00000;
        chicken_boiled[8][5] = 16'b00000_000000_00000;
        chicken_boiled[8][6] = 16'b11111_101000_00100;
        chicken_boiled[8][7] = 16'b11111_101111_01111;
        chicken_boiled[8][8] = 16'b11111_101111_01111;
        chicken_boiled[8][9] = 16'b11111_101111_01111;
        chicken_boiled[8][10] = 16'b11111_101111_01111;
        chicken_boiled[8][11] = 16'b11111_101111_01111;
        chicken_boiled[8][12] = 16'b11111_101000_00100;
        chicken_boiled[8][13] = 16'b00000_000000_00000;
        chicken_boiled[8][14] = 16'b00000_000110_11111;
        chicken_boiled[9][0] = 16'b00000_000110_11111;
        chicken_boiled[9][1] = 16'b00000_000000_00000;
        chicken_boiled[9][2] = 16'b00000_000000_00000;
        chicken_boiled[9][3] = 16'b00000_000000_00000;
        chicken_boiled[9][4] = 16'b00000_000000_00000;
        chicken_boiled[9][5] = 16'b00000_000000_00000;
        chicken_boiled[9][6] = 16'b11111_101000_00100;
        chicken_boiled[9][7] = 16'b11111_101111_01111;
        chicken_boiled[9][8] = 16'b11111_101111_01111;
        chicken_boiled[9][9] = 16'b11111_101111_01111;
        chicken_boiled[9][10] = 16'b11111_101111_01111;
        chicken_boiled[9][11] = 16'b11111_101111_01111;
        chicken_boiled[9][12] = 16'b11111_101000_00100;
        chicken_boiled[9][13] = 16'b11111_101000_00100;
        chicken_boiled[9][14] = 16'b00000_000110_11111;
        chicken_boiled[10][0] = 16'b00000_000110_11111;
        chicken_boiled[10][1] = 16'b00000_000000_00000;
        chicken_boiled[10][2] = 16'b00000_000000_00000;
        chicken_boiled[10][3] = 16'b00000_000000_00000;
        chicken_boiled[10][4] = 16'b00000_000000_00000;
        chicken_boiled[10][5] = 16'b00000_000000_00000;
        chicken_boiled[10][6] = 16'b11111_101000_00100;
        chicken_boiled[10][7] = 16'b11111_101111_01111;
        chicken_boiled[10][8] = 16'b11111_101111_01111;
        chicken_boiled[10][9] = 16'b11111_101111_01111;
        chicken_boiled[10][10] = 16'b11111_101111_01111;
        chicken_boiled[10][11] = 16'b11111_101111_01111;
        chicken_boiled[10][12] = 16'b11111_101111_01111;
        chicken_boiled[10][13] = 16'b11111_101000_00100;
        chicken_boiled[10][14] = 16'b00000_000110_11111;
        chicken_boiled[11][0] = 16'b00000_000110_11111;
        chicken_boiled[11][1] = 16'b00000_000000_00000;
        chicken_boiled[11][2] = 16'b00000_000000_00000;
        chicken_boiled[11][3] = 16'b00000_000000_00000;
        chicken_boiled[11][4] = 16'b00000_000000_00000;
        chicken_boiled[11][5] = 16'b00000_000000_00000;
        chicken_boiled[11][6] = 16'b00000_000000_00000;
        chicken_boiled[11][7] = 16'b11111_101000_00100;
        chicken_boiled[11][8] = 16'b11111_101111_01111;
        chicken_boiled[11][9] = 16'b11111_101111_01111;
        chicken_boiled[11][10] = 16'b11111_101111_01111;
        chicken_boiled[11][11] = 16'b11111_101111_01111;
        chicken_boiled[11][12] = 16'b11111_101000_00100;
        chicken_boiled[11][13] = 16'b11111_101000_00100;
        chicken_boiled[11][14] = 16'b00000_000110_11111;
        chicken_boiled[12][0] = 16'b00000_000110_11111;
        chicken_boiled[12][1] = 16'b00000_000000_00000;
        chicken_boiled[12][2] = 16'b00000_000000_00000;
        chicken_boiled[12][3] = 16'b00000_000000_00000;
        chicken_boiled[12][4] = 16'b00000_000000_00000;
        chicken_boiled[12][5] = 16'b00000_000000_00000;
        chicken_boiled[12][6] = 16'b00000_000000_00000;
        chicken_boiled[12][7] = 16'b11111_101000_00100;
        chicken_boiled[12][8] = 16'b11111_101000_00100;
        chicken_boiled[12][9] = 16'b11111_101111_01111;
        chicken_boiled[12][10] = 16'b11111_101111_01111;
        chicken_boiled[12][11] = 16'b11111_101111_01111;
        chicken_boiled[12][12] = 16'b11111_101000_00100;
        chicken_boiled[12][13] = 16'b00000_000000_00000;
        chicken_boiled[12][14] = 16'b00000_000110_11111;
        chicken_boiled[13][0] = 16'b00000_000110_11111;
        chicken_boiled[13][1] = 16'b00000_000000_00000;
        chicken_boiled[13][2] = 16'b00000_000000_00000;
        chicken_boiled[13][3] = 16'b00000_000000_00000;
        chicken_boiled[13][4] = 16'b00000_000000_00000;
        chicken_boiled[13][5] = 16'b00000_000000_00000;
        chicken_boiled[13][6] = 16'b00000_000000_00000;
        chicken_boiled[13][7] = 16'b00000_000000_00000;
        chicken_boiled[13][8] = 16'b00000_000000_00000;
        chicken_boiled[13][9] = 16'b11111_101000_00100;
        chicken_boiled[13][10] = 16'b11111_101000_00100;
        chicken_boiled[13][11] = 16'b11111_101000_00100;
        chicken_boiled[13][12] = 16'b00000_000000_00000;
        chicken_boiled[13][13] = 16'b00000_000000_00000;
        chicken_boiled[13][14] = 16'b00000_000110_11111;
        chicken_boiled[14][0] = 16'b00000_000110_11111;
        chicken_boiled[14][1] = 16'b00000_000110_11111;
        chicken_boiled[14][2] = 16'b00000_000110_11111;
        chicken_boiled[14][3] = 16'b00000_000110_11111;
        chicken_boiled[14][4] = 16'b00000_000110_11111;
        chicken_boiled[14][5] = 16'b00000_000110_11111;
        chicken_boiled[14][6] = 16'b00000_000110_11111;
        chicken_boiled[14][7] = 16'b00000_000110_11111;
        chicken_boiled[14][8] = 16'b00000_000110_11111;
        chicken_boiled[14][9] = 16'b00000_000110_11111;
        chicken_boiled[14][10] = 16'b00000_000110_11111;
        chicken_boiled[14][11] = 16'b00000_000110_11111;
        chicken_boiled[14][12] = 16'b00000_000110_11111;
        chicken_boiled[14][13] = 16'b00000_000110_11111;
        chicken_boiled[14][14] = 16'b00000_000110_11111;


        chicken_chopped[0][0] = 16'b00000_111111_00001;
        chicken_chopped[0][1] = 16'b00000_111111_00001;
        chicken_chopped[0][2] = 16'b00000_111111_00001;
        chicken_chopped[0][3] = 16'b00000_111111_00001;
        chicken_chopped[0][4] = 16'b00000_111111_00001;
        chicken_chopped[0][5] = 16'b00000_111111_00001;
        chicken_chopped[0][6] = 16'b00000_111111_00001;
        chicken_chopped[0][7] = 16'b00000_111111_00001;
        chicken_chopped[0][8] = 16'b00000_111111_00001;
        chicken_chopped[0][9] = 16'b00000_111111_00001;
        chicken_chopped[0][10] = 16'b00000_111111_00001;
        chicken_chopped[0][11] = 16'b00000_111111_00001;
        chicken_chopped[0][12] = 16'b00000_111111_00001;
        chicken_chopped[0][13] = 16'b00000_111111_00001;
        chicken_chopped[0][14] = 16'b00000_111111_00001;
        chicken_chopped[1][0] = 16'b00000_111111_00001;
        chicken_chopped[1][1] = 16'b11111_111110_11111;
        chicken_chopped[1][2] = 16'b11111_111110_11111;
        chicken_chopped[1][3] = 16'b00000_000000_00000;
        chicken_chopped[1][4] = 16'b00000_000000_00000;
        chicken_chopped[1][5] = 16'b00000_000000_00000;
        chicken_chopped[1][6] = 16'b00000_000000_00000;
        chicken_chopped[1][7] = 16'b00000_000000_00000;
        chicken_chopped[1][8] = 16'b00000_000000_00000;
        chicken_chopped[1][9] = 16'b00000_000000_00000;
        chicken_chopped[1][10] = 16'b00000_000000_00000;
        chicken_chopped[1][11] = 16'b00000_000000_00000;
        chicken_chopped[1][12] = 16'b00000_000000_00000;
        chicken_chopped[1][13] = 16'b00000_000000_00000;
        chicken_chopped[1][14] = 16'b00000_111111_00001;
        chicken_chopped[2][0] = 16'b00000_111111_00001;
        chicken_chopped[2][1] = 16'b11111_111110_11111;
        chicken_chopped[2][2] = 16'b11111_111110_11111;
        chicken_chopped[2][3] = 16'b11111_111110_11111;
        chicken_chopped[2][4] = 16'b00000_000000_00000;
        chicken_chopped[2][5] = 16'b00000_000000_00000;
        chicken_chopped[2][6] = 16'b00000_000000_00000;
        chicken_chopped[2][7] = 16'b00000_000000_00000;
        chicken_chopped[2][8] = 16'b00000_000000_00000;
        chicken_chopped[2][9] = 16'b00000_000000_00000;
        chicken_chopped[2][10] = 16'b00000_000000_00000;
        chicken_chopped[2][11] = 16'b00000_000000_00000;
        chicken_chopped[2][12] = 16'b00000_000000_00000;
        chicken_chopped[2][13] = 16'b00000_000000_00000;
        chicken_chopped[2][14] = 16'b00000_111111_00001;
        chicken_chopped[3][0] = 16'b00000_111111_00001;
        chicken_chopped[3][1] = 16'b00000_000000_00000;
        chicken_chopped[3][2] = 16'b11111_111110_11111;
        chicken_chopped[3][3] = 16'b11111_111110_11111;
        chicken_chopped[3][4] = 16'b11111_111110_11111;
        chicken_chopped[3][5] = 16'b00000_000000_00000;
        chicken_chopped[3][6] = 16'b00000_000000_00000;
        chicken_chopped[3][7] = 16'b00000_000000_00000;
        chicken_chopped[3][8] = 16'b00000_000000_00000;
        chicken_chopped[3][9] = 16'b00000_000000_00000;
        chicken_chopped[3][10] = 16'b00000_000000_00000;
        chicken_chopped[3][11] = 16'b00000_000000_00000;
        chicken_chopped[3][12] = 16'b00000_000000_00000;
        chicken_chopped[3][13] = 16'b00000_000000_00000;
        chicken_chopped[3][14] = 16'b00000_111111_00001;
        chicken_chopped[4][0] = 16'b00000_111111_00001;
        chicken_chopped[4][1] = 16'b00000_000000_00000;
        chicken_chopped[4][2] = 16'b00000_000000_00000;
        chicken_chopped[4][3] = 16'b11111_111110_11111;
        chicken_chopped[4][4] = 16'b11111_101000_00100;
        chicken_chopped[4][5] = 16'b11111_101000_00100;
        chicken_chopped[4][6] = 16'b11111_101000_00100;
        chicken_chopped[4][7] = 16'b00000_000000_00000;
        chicken_chopped[4][8] = 16'b00000_000000_00000;
        chicken_chopped[4][9] = 16'b00000_000000_00000;
        chicken_chopped[4][10] = 16'b00000_000000_00000;
        chicken_chopped[4][11] = 16'b00000_000000_00000;
        chicken_chopped[4][12] = 16'b00000_000000_00000;
        chicken_chopped[4][13] = 16'b00000_000000_00000;
        chicken_chopped[4][14] = 16'b00000_111111_00001;
        chicken_chopped[5][0] = 16'b00000_111111_00001;
        chicken_chopped[5][1] = 16'b00000_000000_00000;
        chicken_chopped[5][2] = 16'b00000_000000_00000;
        chicken_chopped[5][3] = 16'b00000_000000_00000;
        chicken_chopped[5][4] = 16'b11111_101000_00100;
        chicken_chopped[5][5] = 16'b11111_101111_01111;
        chicken_chopped[5][6] = 16'b11111_101111_01111;
        chicken_chopped[5][7] = 16'b11111_101000_00100;
        chicken_chopped[5][8] = 16'b11111_101000_00100;
        chicken_chopped[5][9] = 16'b00000_000000_00000;
        chicken_chopped[5][10] = 16'b00000_000000_00000;
        chicken_chopped[5][11] = 16'b00000_000000_00000;
        chicken_chopped[5][12] = 16'b00000_000000_00000;
        chicken_chopped[5][13] = 16'b00000_000000_00000;
        chicken_chopped[5][14] = 16'b00000_111111_00001;
        chicken_chopped[6][0] = 16'b00000_111111_00001;
        chicken_chopped[6][1] = 16'b00000_000000_00000;
        chicken_chopped[6][2] = 16'b00000_000000_00000;
        chicken_chopped[6][3] = 16'b00000_000000_00000;
        chicken_chopped[6][4] = 16'b00000_000000_00000;
        chicken_chopped[6][5] = 16'b11111_101000_00100;
        chicken_chopped[6][6] = 16'b11111_101111_01111;
        chicken_chopped[6][7] = 16'b11111_101111_01111;
        chicken_chopped[6][8] = 16'b11111_101111_01111;
        chicken_chopped[6][9] = 16'b11111_101000_00100;
        chicken_chopped[6][10] = 16'b11111_101000_00100;
        chicken_chopped[6][11] = 16'b11111_101000_00100;
        chicken_chopped[6][12] = 16'b00000_000000_00000;
        chicken_chopped[6][13] = 16'b00000_000000_00000;
        chicken_chopped[6][14] = 16'b00000_111111_00001;
        chicken_chopped[7][0] = 16'b00000_111111_00001;
        chicken_chopped[7][1] = 16'b00000_000000_00000;
        chicken_chopped[7][2] = 16'b00000_000000_00000;
        chicken_chopped[7][3] = 16'b00000_000000_00000;
        chicken_chopped[7][4] = 16'b00000_000000_00000;
        chicken_chopped[7][5] = 16'b11111_101000_00100;
        chicken_chopped[7][6] = 16'b11111_101111_01111;
        chicken_chopped[7][7] = 16'b11111_101111_01111;
        chicken_chopped[7][8] = 16'b11111_101111_01111;
        chicken_chopped[7][9] = 16'b11111_101111_01111;
        chicken_chopped[7][10] = 16'b11111_101111_01111;
        chicken_chopped[7][11] = 16'b11111_101000_00100;
        chicken_chopped[7][12] = 16'b11111_101000_00100;
        chicken_chopped[7][13] = 16'b00000_000000_00000;
        chicken_chopped[7][14] = 16'b00000_111111_00001;
        chicken_chopped[8][0] = 16'b00000_111111_00001;
        chicken_chopped[8][1] = 16'b00000_000000_00000;
        chicken_chopped[8][2] = 16'b00000_000000_00000;
        chicken_chopped[8][3] = 16'b00000_000000_00000;
        chicken_chopped[8][4] = 16'b00000_000000_00000;
        chicken_chopped[8][5] = 16'b00000_000000_00000;
        chicken_chopped[8][6] = 16'b11111_101000_00100;
        chicken_chopped[8][7] = 16'b11111_101111_01111;
        chicken_chopped[8][8] = 16'b11111_101111_01111;
        chicken_chopped[8][9] = 16'b11111_101111_01111;
        chicken_chopped[8][10] = 16'b11111_101111_01111;
        chicken_chopped[8][11] = 16'b11111_101111_01111;
        chicken_chopped[8][12] = 16'b11111_101000_00100;
        chicken_chopped[8][13] = 16'b00000_000000_00000;
        chicken_chopped[8][14] = 16'b00000_111111_00001;
        chicken_chopped[9][0] = 16'b00000_111111_00001;
        chicken_chopped[9][1] = 16'b00000_000000_00000;
        chicken_chopped[9][2] = 16'b00000_000000_00000;
        chicken_chopped[9][3] = 16'b00000_000000_00000;
        chicken_chopped[9][4] = 16'b00000_000000_00000;
        chicken_chopped[9][5] = 16'b00000_000000_00000;
        chicken_chopped[9][6] = 16'b11111_101000_00100;
        chicken_chopped[9][7] = 16'b11111_101111_01111;
        chicken_chopped[9][8] = 16'b11111_101111_01111;
        chicken_chopped[9][9] = 16'b11111_101111_01111;
        chicken_chopped[9][10] = 16'b11111_101111_01111;
        chicken_chopped[9][11] = 16'b11111_101111_01111;
        chicken_chopped[9][12] = 16'b11111_101000_00100;
        chicken_chopped[9][13] = 16'b11111_101000_00100;
        chicken_chopped[9][14] = 16'b00000_111111_00001;
        chicken_chopped[10][0] = 16'b00000_111111_00001;
        chicken_chopped[10][1] = 16'b00000_000000_00000;
        chicken_chopped[10][2] = 16'b00000_000000_00000;
        chicken_chopped[10][3] = 16'b00000_000000_00000;
        chicken_chopped[10][4] = 16'b00000_000000_00000;
        chicken_chopped[10][5] = 16'b00000_000000_00000;
        chicken_chopped[10][6] = 16'b11111_101000_00100;
        chicken_chopped[10][7] = 16'b11111_101111_01111;
        chicken_chopped[10][8] = 16'b11111_101111_01111;
        chicken_chopped[10][9] = 16'b11111_101111_01111;
        chicken_chopped[10][10] = 16'b11111_101111_01111;
        chicken_chopped[10][11] = 16'b11111_101111_01111;
        chicken_chopped[10][12] = 16'b11111_101111_01111;
        chicken_chopped[10][13] = 16'b11111_101000_00100;
        chicken_chopped[10][14] = 16'b00000_111111_00001;
        chicken_chopped[11][0] = 16'b00000_111111_00001;
        chicken_chopped[11][1] = 16'b00000_000000_00000;
        chicken_chopped[11][2] = 16'b00000_000000_00000;
        chicken_chopped[11][3] = 16'b00000_000000_00000;
        chicken_chopped[11][4] = 16'b00000_000000_00000;
        chicken_chopped[11][5] = 16'b00000_000000_00000;
        chicken_chopped[11][6] = 16'b00000_000000_00000;
        chicken_chopped[11][7] = 16'b11111_101000_00100;
        chicken_chopped[11][8] = 16'b11111_101111_01111;
        chicken_chopped[11][9] = 16'b11111_101111_01111;
        chicken_chopped[11][10] = 16'b11111_101111_01111;
        chicken_chopped[11][11] = 16'b11111_101111_01111;
        chicken_chopped[11][12] = 16'b11111_101000_00100;
        chicken_chopped[11][13] = 16'b11111_101000_00100;
        chicken_chopped[11][14] = 16'b00000_111111_00001;
        chicken_chopped[12][0] = 16'b00000_111111_00001;
        chicken_chopped[12][1] = 16'b00000_000000_00000;
        chicken_chopped[12][2] = 16'b00000_000000_00000;
        chicken_chopped[12][3] = 16'b00000_000000_00000;
        chicken_chopped[12][4] = 16'b00000_000000_00000;
        chicken_chopped[12][5] = 16'b00000_000000_00000;
        chicken_chopped[12][6] = 16'b00000_000000_00000;
        chicken_chopped[12][7] = 16'b11111_101000_00100;
        chicken_chopped[12][8] = 16'b11111_101000_00100;
        chicken_chopped[12][9] = 16'b11111_101111_01111;
        chicken_chopped[12][10] = 16'b11111_101111_01111;
        chicken_chopped[12][11] = 16'b11111_101111_01111;
        chicken_chopped[12][12] = 16'b11111_101000_00100;
        chicken_chopped[12][13] = 16'b00000_000000_00000;
        chicken_chopped[12][14] = 16'b00000_111111_00001;
        chicken_chopped[13][0] = 16'b00000_111111_00001;
        chicken_chopped[13][1] = 16'b00000_000000_00000;
        chicken_chopped[13][2] = 16'b00000_000000_00000;
        chicken_chopped[13][3] = 16'b00000_000000_00000;
        chicken_chopped[13][4] = 16'b00000_000000_00000;
        chicken_chopped[13][5] = 16'b00000_000000_00000;
        chicken_chopped[13][6] = 16'b00000_000000_00000;
        chicken_chopped[13][7] = 16'b00000_000000_00000;
        chicken_chopped[13][8] = 16'b00000_000000_00000;
        chicken_chopped[13][9] = 16'b11111_101000_00100;
        chicken_chopped[13][10] = 16'b11111_101000_00100;
        chicken_chopped[13][11] = 16'b11111_101000_00100;
        chicken_chopped[13][12] = 16'b00000_000000_00000;
        chicken_chopped[13][13] = 16'b00000_000000_00000;
        chicken_chopped[13][14] = 16'b00000_111111_00001;
        chicken_chopped[14][0] = 16'b00000_111111_00001;
        chicken_chopped[14][1] = 16'b00000_111111_00001;
        chicken_chopped[14][2] = 16'b00000_111111_00001;
        chicken_chopped[14][3] = 16'b00000_111111_00001;
        chicken_chopped[14][4] = 16'b00000_111111_00001;
        chicken_chopped[14][5] = 16'b00000_111111_00001;
        chicken_chopped[14][6] = 16'b00000_111111_00001;
        chicken_chopped[14][7] = 16'b00000_111111_00001;
        chicken_chopped[14][8] = 16'b00000_111111_00001;
        chicken_chopped[14][9] = 16'b00000_111111_00001;
        chicken_chopped[14][10] = 16'b00000_111111_00001;
        chicken_chopped[14][11] = 16'b00000_111111_00001;
        chicken_chopped[14][12] = 16'b00000_111111_00001;
        chicken_chopped[14][13] = 16'b00000_111111_00001;
        chicken_chopped[14][14] = 16'b00000_111111_00001;


        chicken_raw[0][0] = 16'b11111_101111_01111;
        chicken_raw[0][1] = 16'b11111_101111_01111;
        chicken_raw[0][2] = 16'b11111_101111_01111;
        chicken_raw[0][3] = 16'b11111_101111_01111;
        chicken_raw[0][4] = 16'b11111_101111_01111;
        chicken_raw[0][5] = 16'b11111_101111_01111;
        chicken_raw[0][6] = 16'b11111_101111_01111;
        chicken_raw[0][7] = 16'b11111_101111_01111;
        chicken_raw[0][8] = 16'b11111_101111_01111;
        chicken_raw[0][9] = 16'b11111_101111_01111;
        chicken_raw[0][10] = 16'b11111_101111_01111;
        chicken_raw[0][11] = 16'b11111_101111_01111;
        chicken_raw[0][12] = 16'b11111_101111_01111;
        chicken_raw[0][13] = 16'b11111_101111_01111;
        chicken_raw[0][14] = 16'b11111_101111_01111;
        chicken_raw[1][0] = 16'b11111_101111_01111;
        chicken_raw[1][1] = 16'b11111_111110_11111;
        chicken_raw[1][2] = 16'b11111_111110_11111;
        chicken_raw[1][3] = 16'b00000_000000_00000;
        chicken_raw[1][4] = 16'b00000_000000_00000;
        chicken_raw[1][5] = 16'b00000_000000_00000;
        chicken_raw[1][6] = 16'b00000_000000_00000;
        chicken_raw[1][7] = 16'b00000_000000_00000;
        chicken_raw[1][8] = 16'b00000_000000_00000;
        chicken_raw[1][9] = 16'b00000_000000_00000;
        chicken_raw[1][10] = 16'b00000_000000_00000;
        chicken_raw[1][11] = 16'b00000_000000_00000;
        chicken_raw[1][12] = 16'b00000_000000_00000;
        chicken_raw[1][13] = 16'b00000_000000_00000;
        chicken_raw[1][14] = 16'b11111_101111_01111;
        chicken_raw[2][0] = 16'b11111_101111_01111;
        chicken_raw[2][1] = 16'b11111_111110_11111;
        chicken_raw[2][2] = 16'b11111_111110_11111;
        chicken_raw[2][3] = 16'b11111_111110_11111;
        chicken_raw[2][4] = 16'b00000_000000_00000;
        chicken_raw[2][5] = 16'b00000_000000_00000;
        chicken_raw[2][6] = 16'b00000_000000_00000;
        chicken_raw[2][7] = 16'b00000_000000_00000;
        chicken_raw[2][8] = 16'b00000_000000_00000;
        chicken_raw[2][9] = 16'b00000_000000_00000;
        chicken_raw[2][10] = 16'b00000_000000_00000;
        chicken_raw[2][11] = 16'b00000_000000_00000;
        chicken_raw[2][12] = 16'b00000_000000_00000;
        chicken_raw[2][13] = 16'b00000_000000_00000;
        chicken_raw[2][14] = 16'b11111_101111_01111;
        chicken_raw[3][0] = 16'b11111_101111_01111;
        chicken_raw[3][1] = 16'b00000_000000_00000;
        chicken_raw[3][2] = 16'b11111_111110_11111;
        chicken_raw[3][3] = 16'b11111_111110_11111;
        chicken_raw[3][4] = 16'b11111_111110_11111;
        chicken_raw[3][5] = 16'b00000_000000_00000;
        chicken_raw[3][6] = 16'b00000_000000_00000;
        chicken_raw[3][7] = 16'b00000_000000_00000;
        chicken_raw[3][8] = 16'b00000_000000_00000;
        chicken_raw[3][9] = 16'b00000_000000_00000;
        chicken_raw[3][10] = 16'b00000_000000_00000;
        chicken_raw[3][11] = 16'b00000_000000_00000;
        chicken_raw[3][12] = 16'b00000_000000_00000;
        chicken_raw[3][13] = 16'b00000_000000_00000;
        chicken_raw[3][14] = 16'b11111_101111_01111;
        chicken_raw[4][0] = 16'b11111_101111_01111;
        chicken_raw[4][1] = 16'b00000_000000_00000;
        chicken_raw[4][2] = 16'b00000_000000_00000;
        chicken_raw[4][3] = 16'b11111_111110_11111;
        chicken_raw[4][4] = 16'b11111_101000_00100;
        chicken_raw[4][5] = 16'b11111_101000_00100;
        chicken_raw[4][6] = 16'b11111_101000_00100;
        chicken_raw[4][7] = 16'b00000_000000_00000;
        chicken_raw[4][8] = 16'b00000_000000_00000;
        chicken_raw[4][9] = 16'b00000_000000_00000;
        chicken_raw[4][10] = 16'b00000_000000_00000;
        chicken_raw[4][11] = 16'b00000_000000_00000;
        chicken_raw[4][12] = 16'b00000_000000_00000;
        chicken_raw[4][13] = 16'b00000_000000_00000;
        chicken_raw[4][14] = 16'b11111_101111_01111;
        chicken_raw[5][0] = 16'b11111_101111_01111;
        chicken_raw[5][1] = 16'b00000_000000_00000;
        chicken_raw[5][2] = 16'b00000_000000_00000;
        chicken_raw[5][3] = 16'b00000_000000_00000;
        chicken_raw[5][4] = 16'b11111_101000_00100;
        chicken_raw[5][5] = 16'b11111_101111_01111;
        chicken_raw[5][6] = 16'b11111_101111_01111;
        chicken_raw[5][7] = 16'b11111_101000_00100;
        chicken_raw[5][8] = 16'b11111_101000_00100;
        chicken_raw[5][9] = 16'b00000_000000_00000;
        chicken_raw[5][10] = 16'b00000_000000_00000;
        chicken_raw[5][11] = 16'b00000_000000_00000;
        chicken_raw[5][12] = 16'b00000_000000_00000;
        chicken_raw[5][13] = 16'b00000_000000_00000;
        chicken_raw[5][14] = 16'b11111_101111_01111;
        chicken_raw[6][0] = 16'b11111_101111_01111;
        chicken_raw[6][1] = 16'b00000_000000_00000;
        chicken_raw[6][2] = 16'b00000_000000_00000;
        chicken_raw[6][3] = 16'b00000_000000_00000;
        chicken_raw[6][4] = 16'b00000_000000_00000;
        chicken_raw[6][5] = 16'b11111_101000_00100;
        chicken_raw[6][6] = 16'b11111_101111_01111;
        chicken_raw[6][7] = 16'b11111_101111_01111;
        chicken_raw[6][8] = 16'b11111_101111_01111;
        chicken_raw[6][9] = 16'b11111_101000_00100;
        chicken_raw[6][10] = 16'b11111_101000_00100;
        chicken_raw[6][11] = 16'b11111_101000_00100;
        chicken_raw[6][12] = 16'b00000_000000_00000;
        chicken_raw[6][13] = 16'b00000_000000_00000;
        chicken_raw[6][14] = 16'b11111_101111_01111;
        chicken_raw[7][0] = 16'b11111_101111_01111;
        chicken_raw[7][1] = 16'b00000_000000_00000;
        chicken_raw[7][2] = 16'b00000_000000_00000;
        chicken_raw[7][3] = 16'b00000_000000_00000;
        chicken_raw[7][4] = 16'b00000_000000_00000;
        chicken_raw[7][5] = 16'b11111_101000_00100;
        chicken_raw[7][6] = 16'b11111_101111_01111;
        chicken_raw[7][7] = 16'b11111_101111_01111;
        chicken_raw[7][8] = 16'b11111_101111_01111;
        chicken_raw[7][9] = 16'b11111_101111_01111;
        chicken_raw[7][10] = 16'b11111_101111_01111;
        chicken_raw[7][11] = 16'b11111_101000_00100;
        chicken_raw[7][12] = 16'b11111_101000_00100;
        chicken_raw[7][13] = 16'b00000_000000_00000;
        chicken_raw[7][14] = 16'b11111_101111_01111;
        chicken_raw[8][0] = 16'b11111_101111_01111;
        chicken_raw[8][1] = 16'b00000_000000_00000;
        chicken_raw[8][2] = 16'b00000_000000_00000;
        chicken_raw[8][3] = 16'b00000_000000_00000;
        chicken_raw[8][4] = 16'b00000_000000_00000;
        chicken_raw[8][5] = 16'b00000_000000_00000;
        chicken_raw[8][6] = 16'b11111_101000_00100;
        chicken_raw[8][7] = 16'b11111_101111_01111;
        chicken_raw[8][8] = 16'b11111_101111_01111;
        chicken_raw[8][9] = 16'b11111_101111_01111;
        chicken_raw[8][10] = 16'b11111_101111_01111;
        chicken_raw[8][11] = 16'b11111_101111_01111;
        chicken_raw[8][12] = 16'b11111_101000_00100;
        chicken_raw[8][13] = 16'b00000_000000_00000;
        chicken_raw[8][14] = 16'b11111_101111_01111;
        chicken_raw[9][0] = 16'b11111_101111_01111;
        chicken_raw[9][1] = 16'b00000_000000_00000;
        chicken_raw[9][2] = 16'b00000_000000_00000;
        chicken_raw[9][3] = 16'b00000_000000_00000;
        chicken_raw[9][4] = 16'b00000_000000_00000;
        chicken_raw[9][5] = 16'b00000_000000_00000;
        chicken_raw[9][6] = 16'b11111_101000_00100;
        chicken_raw[9][7] = 16'b11111_101111_01111;
        chicken_raw[9][8] = 16'b11111_101111_01111;
        chicken_raw[9][9] = 16'b11111_101111_01111;
        chicken_raw[9][10] = 16'b11111_101111_01111;
        chicken_raw[9][11] = 16'b11111_101111_01111;
        chicken_raw[9][12] = 16'b11111_101000_00100;
        chicken_raw[9][13] = 16'b11111_101000_00100;
        chicken_raw[9][14] = 16'b11111_101111_01111;
        chicken_raw[10][0] = 16'b11111_101111_01111;
        chicken_raw[10][1] = 16'b00000_000000_00000;
        chicken_raw[10][2] = 16'b00000_000000_00000;
        chicken_raw[10][3] = 16'b00000_000000_00000;
        chicken_raw[10][4] = 16'b00000_000000_00000;
        chicken_raw[10][5] = 16'b00000_000000_00000;
        chicken_raw[10][6] = 16'b11111_101000_00100;
        chicken_raw[10][7] = 16'b11111_101111_01111;
        chicken_raw[10][8] = 16'b11111_101111_01111;
        chicken_raw[10][9] = 16'b11111_101111_01111;
        chicken_raw[10][10] = 16'b11111_101111_01111;
        chicken_raw[10][11] = 16'b11111_101111_01111;
        chicken_raw[10][12] = 16'b11111_101111_01111;
        chicken_raw[10][13] = 16'b11111_101000_00100;
        chicken_raw[10][14] = 16'b11111_101111_01111;
        chicken_raw[11][0] = 16'b11111_101111_01111;
        chicken_raw[11][1] = 16'b00000_000000_00000;
        chicken_raw[11][2] = 16'b00000_000000_00000;
        chicken_raw[11][3] = 16'b00000_000000_00000;
        chicken_raw[11][4] = 16'b00000_000000_00000;
        chicken_raw[11][5] = 16'b00000_000000_00000;
        chicken_raw[11][6] = 16'b00000_000000_00000;
        chicken_raw[11][7] = 16'b11111_101000_00100;
        chicken_raw[11][8] = 16'b11111_101111_01111;
        chicken_raw[11][9] = 16'b11111_101111_01111;
        chicken_raw[11][10] = 16'b11111_101111_01111;
        chicken_raw[11][11] = 16'b11111_101111_01111;
        chicken_raw[11][12] = 16'b11111_101000_00100;
        chicken_raw[11][13] = 16'b11111_101000_00100;
        chicken_raw[11][14] = 16'b11111_101111_01111;
        chicken_raw[12][0] = 16'b11111_101111_01111;
        chicken_raw[12][1] = 16'b00000_000000_00000;
        chicken_raw[12][2] = 16'b00000_000000_00000;
        chicken_raw[12][3] = 16'b00000_000000_00000;
        chicken_raw[12][4] = 16'b00000_000000_00000;
        chicken_raw[12][5] = 16'b00000_000000_00000;
        chicken_raw[12][6] = 16'b00000_000000_00000;
        chicken_raw[12][7] = 16'b11111_101000_00100;
        chicken_raw[12][8] = 16'b11111_101000_00100;
        chicken_raw[12][9] = 16'b11111_101111_01111;
        chicken_raw[12][10] = 16'b11111_101111_01111;
        chicken_raw[12][11] = 16'b11111_101111_01111;
        chicken_raw[12][12] = 16'b11111_101000_00100;
        chicken_raw[12][13] = 16'b00000_000000_00000;
        chicken_raw[12][14] = 16'b11111_101111_01111;
        chicken_raw[13][0] = 16'b11111_101111_01111;
        chicken_raw[13][1] = 16'b00000_000000_00000;
        chicken_raw[13][2] = 16'b00000_000000_00000;
        chicken_raw[13][3] = 16'b00000_000000_00000;
        chicken_raw[13][4] = 16'b00000_000000_00000;
        chicken_raw[13][5] = 16'b00000_000000_00000;
        chicken_raw[13][6] = 16'b00000_000000_00000;
        chicken_raw[13][7] = 16'b00000_000000_00000;
        chicken_raw[13][8] = 16'b00000_000000_00000;
        chicken_raw[13][9] = 16'b11111_101000_00100;
        chicken_raw[13][10] = 16'b11111_101000_00100;
        chicken_raw[13][11] = 16'b11111_101000_00100;
        chicken_raw[13][12] = 16'b00000_000000_00000;
        chicken_raw[13][13] = 16'b00000_000000_00000;
        chicken_raw[13][14] = 16'b11111_101111_01111;
        chicken_raw[14][0] = 16'b11111_101111_01111;
        chicken_raw[14][1] = 16'b11111_101111_01111;
        chicken_raw[14][2] = 16'b11111_101111_01111;
        chicken_raw[14][3] = 16'b11111_101111_01111;
        chicken_raw[14][4] = 16'b11111_101111_01111;
        chicken_raw[14][5] = 16'b11111_101111_01111;
        chicken_raw[14][6] = 16'b11111_101111_01111;
        chicken_raw[14][7] = 16'b11111_101111_01111;
        chicken_raw[14][8] = 16'b11111_101111_01111;
        chicken_raw[14][9] = 16'b11111_101111_01111;
        chicken_raw[14][10] = 16'b11111_101111_01111;
        chicken_raw[14][11] = 16'b11111_101111_01111;
        chicken_raw[14][12] = 16'b11111_101111_01111;
        chicken_raw[14][13] = 16'b11111_101111_01111;
        chicken_raw[14][14] = 16'b11111_101111_01111;


        onion_boiled_chopped[0][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][1] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][2] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][3] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][4] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][5] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][6] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][7] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][8] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][9] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][10] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][11] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][12] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][13] = 16'b10101_011000_00000;
        onion_boiled_chopped[0][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[1][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[1][1] = 16'b00000_000000_00000;
        onion_boiled_chopped[1][2] = 16'b00000_000000_00000;
        onion_boiled_chopped[1][3] = 16'b10100_000000_11111;
        onion_boiled_chopped[1][4] = 16'b10100_000000_11111;
        onion_boiled_chopped[1][5] = 16'b10100_000000_11111;
        onion_boiled_chopped[1][6] = 16'b10100_000000_11111;
        onion_boiled_chopped[1][7] = 16'b10100_000000_11111;
        onion_boiled_chopped[1][8] = 16'b10100_000000_11111;
        onion_boiled_chopped[1][9] = 16'b10100_000000_11111;
        onion_boiled_chopped[1][10] = 16'b10100_000000_11111;
        onion_boiled_chopped[1][11] = 16'b00000_000000_00000;
        onion_boiled_chopped[1][12] = 16'b00000_000000_00000;
        onion_boiled_chopped[1][13] = 16'b00000_000000_00000;
        onion_boiled_chopped[1][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[2][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[2][1] = 16'b00000_000000_00000;
        onion_boiled_chopped[2][2] = 16'b10100_000000_11111;
        onion_boiled_chopped[2][3] = 16'b10100_000000_11111;
        onion_boiled_chopped[2][4] = 16'b11001_100101_11111;
        onion_boiled_chopped[2][5] = 16'b11001_100101_11111;
        onion_boiled_chopped[2][6] = 16'b11001_100101_11111;
        onion_boiled_chopped[2][7] = 16'b11001_100101_11111;
        onion_boiled_chopped[2][8] = 16'b11001_100101_11111;
        onion_boiled_chopped[2][9] = 16'b11001_100101_11111;
        onion_boiled_chopped[2][10] = 16'b11001_100101_11111;
        onion_boiled_chopped[2][11] = 16'b11001_100101_11111;
        onion_boiled_chopped[2][12] = 16'b10100_000000_11111;
        onion_boiled_chopped[2][13] = 16'b00000_000000_00000;
        onion_boiled_chopped[2][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[3][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[3][1] = 16'b10100_000000_11111;
        onion_boiled_chopped[3][2] = 16'b10100_000000_11111;
        onion_boiled_chopped[3][3] = 16'b11001_100101_11111;
        onion_boiled_chopped[3][4] = 16'b10100_000000_11111;
        onion_boiled_chopped[3][5] = 16'b10100_000000_11111;
        onion_boiled_chopped[3][6] = 16'b10100_000000_11111;
        onion_boiled_chopped[3][7] = 16'b10100_000000_11111;
        onion_boiled_chopped[3][8] = 16'b10100_000000_11111;
        onion_boiled_chopped[3][9] = 16'b10100_000000_11111;
        onion_boiled_chopped[3][10] = 16'b10100_000000_11111;
        onion_boiled_chopped[3][11] = 16'b11001_100101_11111;
        onion_boiled_chopped[3][12] = 16'b10100_000000_11111;
        onion_boiled_chopped[3][13] = 16'b00000_000000_00000;
        onion_boiled_chopped[3][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[4][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[4][1] = 16'b10100_000000_11111;
        onion_boiled_chopped[4][2] = 16'b11001_100101_11111;
        onion_boiled_chopped[4][3] = 16'b10100_000000_11111;
        onion_boiled_chopped[4][4] = 16'b10100_000000_11111;
        onion_boiled_chopped[4][5] = 16'b11001_100101_11111;
        onion_boiled_chopped[4][6] = 16'b11001_100101_11111;
        onion_boiled_chopped[4][7] = 16'b11001_100101_11111;
        onion_boiled_chopped[4][8] = 16'b11001_100101_11111;
        onion_boiled_chopped[4][9] = 16'b11001_100101_11111;
        onion_boiled_chopped[4][10] = 16'b10100_000000_11111;
        onion_boiled_chopped[4][11] = 16'b10100_000000_11111;
        onion_boiled_chopped[4][12] = 16'b11001_100101_11111;
        onion_boiled_chopped[4][13] = 16'b10100_000000_11111;
        onion_boiled_chopped[4][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[5][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[5][1] = 16'b10100_000000_11111;
        onion_boiled_chopped[5][2] = 16'b11001_100101_11111;
        onion_boiled_chopped[5][3] = 16'b10100_000000_11111;
        onion_boiled_chopped[5][4] = 16'b11001_100101_11111;
        onion_boiled_chopped[5][5] = 16'b10100_000000_11111;
        onion_boiled_chopped[5][6] = 16'b10100_000000_11111;
        onion_boiled_chopped[5][7] = 16'b10100_000000_11111;
        onion_boiled_chopped[5][8] = 16'b10100_000000_11111;
        onion_boiled_chopped[5][9] = 16'b10100_000000_11111;
        onion_boiled_chopped[5][10] = 16'b11001_100101_11111;
        onion_boiled_chopped[5][11] = 16'b10100_000000_11111;
        onion_boiled_chopped[5][12] = 16'b11001_100101_11111;
        onion_boiled_chopped[5][13] = 16'b10100_000000_11111;
        onion_boiled_chopped[5][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[6][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[6][1] = 16'b10100_000000_11111;
        onion_boiled_chopped[6][2] = 16'b11001_100101_11111;
        onion_boiled_chopped[6][3] = 16'b10100_000000_11111;
        onion_boiled_chopped[6][4] = 16'b11001_100101_11111;
        onion_boiled_chopped[6][5] = 16'b10100_000000_11111;
        onion_boiled_chopped[6][6] = 16'b10100_000000_11111;
        onion_boiled_chopped[6][7] = 16'b11001_100101_11111;
        onion_boiled_chopped[6][8] = 16'b10100_000000_11111;
        onion_boiled_chopped[6][9] = 16'b10100_000000_11111;
        onion_boiled_chopped[6][10] = 16'b11001_100101_11111;
        onion_boiled_chopped[6][11] = 16'b10100_000000_11111;
        onion_boiled_chopped[6][12] = 16'b11001_100101_11111;
        onion_boiled_chopped[6][13] = 16'b10100_000000_11111;
        onion_boiled_chopped[6][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[7][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[7][1] = 16'b00000_000000_00000;
        onion_boiled_chopped[7][2] = 16'b11001_100101_11111;
        onion_boiled_chopped[7][3] = 16'b10100_000000_11111;
        onion_boiled_chopped[7][4] = 16'b10100_000000_11111;
        onion_boiled_chopped[7][5] = 16'b11001_100101_11111;
        onion_boiled_chopped[7][6] = 16'b10100_000000_11111;
        onion_boiled_chopped[7][7] = 16'b10100_000000_11111;
        onion_boiled_chopped[7][8] = 16'b11001_100101_11111;
        onion_boiled_chopped[7][9] = 16'b10100_000000_11111;
        onion_boiled_chopped[7][10] = 16'b11001_100101_11111;
        onion_boiled_chopped[7][11] = 16'b10100_000000_11111;
        onion_boiled_chopped[7][12] = 16'b11001_100101_11111;
        onion_boiled_chopped[7][13] = 16'b10100_000000_11111;
        onion_boiled_chopped[7][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[8][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[8][1] = 16'b00000_000000_00000;
        onion_boiled_chopped[8][2] = 16'b10100_000000_11111;
        onion_boiled_chopped[8][3] = 16'b11001_100101_11111;
        onion_boiled_chopped[8][4] = 16'b10100_000000_11111;
        onion_boiled_chopped[8][5] = 16'b10100_000000_11111;
        onion_boiled_chopped[8][6] = 16'b11001_100101_11111;
        onion_boiled_chopped[8][7] = 16'b10100_000000_11111;
        onion_boiled_chopped[8][8] = 16'b10100_000000_11111;
        onion_boiled_chopped[8][9] = 16'b11001_100101_11111;
        onion_boiled_chopped[8][10] = 16'b10100_000000_11111;
        onion_boiled_chopped[8][11] = 16'b10100_000000_11111;
        onion_boiled_chopped[8][12] = 16'b11001_100101_11111;
        onion_boiled_chopped[8][13] = 16'b10100_000000_11111;
        onion_boiled_chopped[8][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[9][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[9][1] = 16'b00000_000000_00000;
        onion_boiled_chopped[9][2] = 16'b00000_000000_00000;
        onion_boiled_chopped[9][3] = 16'b10100_000000_11111;
        onion_boiled_chopped[9][4] = 16'b11001_100101_11111;
        onion_boiled_chopped[9][5] = 16'b10100_000000_11111;
        onion_boiled_chopped[9][6] = 16'b10100_000000_11111;
        onion_boiled_chopped[9][7] = 16'b11001_100101_11111;
        onion_boiled_chopped[9][8] = 16'b11001_100101_11111;
        onion_boiled_chopped[9][9] = 16'b10100_000000_11111;
        onion_boiled_chopped[9][10] = 16'b10100_000000_11111;
        onion_boiled_chopped[9][11] = 16'b11001_100101_11111;
        onion_boiled_chopped[9][12] = 16'b10100_000000_11111;
        onion_boiled_chopped[9][13] = 16'b00000_000000_00000;
        onion_boiled_chopped[9][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[10][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[10][1] = 16'b00000_000000_00000;
        onion_boiled_chopped[10][2] = 16'b00000_000000_00000;
        onion_boiled_chopped[10][3] = 16'b00000_000000_00000;
        onion_boiled_chopped[10][4] = 16'b10100_000000_11111;
        onion_boiled_chopped[10][5] = 16'b11001_100101_11111;
        onion_boiled_chopped[10][6] = 16'b10100_000000_11111;
        onion_boiled_chopped[10][7] = 16'b10100_000000_11111;
        onion_boiled_chopped[10][8] = 16'b10100_000000_11111;
        onion_boiled_chopped[10][9] = 16'b10100_000000_11111;
        onion_boiled_chopped[10][10] = 16'b11001_100101_11111;
        onion_boiled_chopped[10][11] = 16'b10100_000000_11111;
        onion_boiled_chopped[10][12] = 16'b00000_000000_00000;
        onion_boiled_chopped[10][13] = 16'b00000_000000_00000;
        onion_boiled_chopped[10][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[11][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[11][1] = 16'b00000_000000_00000;
        onion_boiled_chopped[11][2] = 16'b00000_000000_00000;
        onion_boiled_chopped[11][3] = 16'b00000_000000_00000;
        onion_boiled_chopped[11][4] = 16'b00000_000000_00000;
        onion_boiled_chopped[11][5] = 16'b10100_000000_11111;
        onion_boiled_chopped[11][6] = 16'b11001_100101_11111;
        onion_boiled_chopped[11][7] = 16'b10100_000000_11111;
        onion_boiled_chopped[11][8] = 16'b10100_000000_11111;
        onion_boiled_chopped[11][9] = 16'b11001_100101_11111;
        onion_boiled_chopped[11][10] = 16'b10100_000000_11111;
        onion_boiled_chopped[11][11] = 16'b00000_000000_00000;
        onion_boiled_chopped[11][12] = 16'b00000_000000_00000;
        onion_boiled_chopped[11][13] = 16'b00000_000000_00000;
        onion_boiled_chopped[11][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[12][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[12][1] = 16'b00000_000000_00000;
        onion_boiled_chopped[12][2] = 16'b00000_000000_00000;
        onion_boiled_chopped[12][3] = 16'b00000_000000_00000;
        onion_boiled_chopped[12][4] = 16'b00000_000000_00000;
        onion_boiled_chopped[12][5] = 16'b00000_000000_00000;
        onion_boiled_chopped[12][6] = 16'b10100_000000_11111;
        onion_boiled_chopped[12][7] = 16'b11001_100101_11111;
        onion_boiled_chopped[12][8] = 16'b11001_100101_11111;
        onion_boiled_chopped[12][9] = 16'b10100_000000_11111;
        onion_boiled_chopped[12][10] = 16'b00000_000000_00000;
        onion_boiled_chopped[12][11] = 16'b00000_000000_00000;
        onion_boiled_chopped[12][12] = 16'b00000_000000_00000;
        onion_boiled_chopped[12][13] = 16'b00000_000000_00000;
        onion_boiled_chopped[12][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[13][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[13][1] = 16'b00000_000000_00000;
        onion_boiled_chopped[13][2] = 16'b00000_000000_00000;
        onion_boiled_chopped[13][3] = 16'b00000_000000_00000;
        onion_boiled_chopped[13][4] = 16'b00000_000000_00000;
        onion_boiled_chopped[13][5] = 16'b00000_000000_00000;
        onion_boiled_chopped[13][6] = 16'b00000_000000_00000;
        onion_boiled_chopped[13][7] = 16'b10100_000000_11111;
        onion_boiled_chopped[13][8] = 16'b00000_000000_00000;
        onion_boiled_chopped[13][9] = 16'b00000_000000_00000;
        onion_boiled_chopped[13][10] = 16'b00000_000000_00000;
        onion_boiled_chopped[13][11] = 16'b00000_000000_00000;
        onion_boiled_chopped[13][12] = 16'b00000_000000_00000;
        onion_boiled_chopped[13][13] = 16'b00000_000000_00000;
        onion_boiled_chopped[13][14] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][0] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][1] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][2] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][3] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][4] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][5] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][6] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][7] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][8] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][9] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][10] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][11] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][12] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][13] = 16'b10101_011000_00000;
        onion_boiled_chopped[14][14] = 16'b10101_011000_00000;


        onion_boiled[0][0] = 16'b00000_000110_11111;
        onion_boiled[0][1] = 16'b00000_000110_11111;
        onion_boiled[0][2] = 16'b00000_000110_11111;
        onion_boiled[0][3] = 16'b00000_000110_11111;
        onion_boiled[0][4] = 16'b00000_000110_11111;
        onion_boiled[0][5] = 16'b00000_000110_11111;
        onion_boiled[0][6] = 16'b00000_000110_11111;
        onion_boiled[0][7] = 16'b00000_000110_11111;
        onion_boiled[0][8] = 16'b00000_000110_11111;
        onion_boiled[0][9] = 16'b00000_000110_11111;
        onion_boiled[0][10] = 16'b00000_000110_11111;
        onion_boiled[0][11] = 16'b00000_000110_11111;
        onion_boiled[0][12] = 16'b00000_000110_11111;
        onion_boiled[0][13] = 16'b00000_000110_11111;
        onion_boiled[0][14] = 16'b00000_000110_11111;
        onion_boiled[1][0] = 16'b00000_000110_11111;
        onion_boiled[1][1] = 16'b00000_000000_00000;
        onion_boiled[1][2] = 16'b00000_000000_00000;
        onion_boiled[1][3] = 16'b10100_000000_11111;
        onion_boiled[1][4] = 16'b10100_000000_11111;
        onion_boiled[1][5] = 16'b10100_000000_11111;
        onion_boiled[1][6] = 16'b10100_000000_11111;
        onion_boiled[1][7] = 16'b10100_000000_11111;
        onion_boiled[1][8] = 16'b10100_000000_11111;
        onion_boiled[1][9] = 16'b10100_000000_11111;
        onion_boiled[1][10] = 16'b10100_000000_11111;
        onion_boiled[1][11] = 16'b00000_000000_00000;
        onion_boiled[1][12] = 16'b00000_000000_00000;
        onion_boiled[1][13] = 16'b00000_000000_00000;
        onion_boiled[1][14] = 16'b00000_000110_11111;
        onion_boiled[2][0] = 16'b00000_000110_11111;
        onion_boiled[2][1] = 16'b00000_000000_00000;
        onion_boiled[2][2] = 16'b10100_000000_11111;
        onion_boiled[2][3] = 16'b10100_000000_11111;
        onion_boiled[2][4] = 16'b11001_100101_11111;
        onion_boiled[2][5] = 16'b11001_100101_11111;
        onion_boiled[2][6] = 16'b11001_100101_11111;
        onion_boiled[2][7] = 16'b11001_100101_11111;
        onion_boiled[2][8] = 16'b11001_100101_11111;
        onion_boiled[2][9] = 16'b11001_100101_11111;
        onion_boiled[2][10] = 16'b11001_100101_11111;
        onion_boiled[2][11] = 16'b11001_100101_11111;
        onion_boiled[2][12] = 16'b10100_000000_11111;
        onion_boiled[2][13] = 16'b00000_000000_00000;
        onion_boiled[2][14] = 16'b00000_000110_11111;
        onion_boiled[3][0] = 16'b00000_000110_11111;
        onion_boiled[3][1] = 16'b10100_000000_11111;
        onion_boiled[3][2] = 16'b10100_000000_11111;
        onion_boiled[3][3] = 16'b11001_100101_11111;
        onion_boiled[3][4] = 16'b10100_000000_11111;
        onion_boiled[3][5] = 16'b10100_000000_11111;
        onion_boiled[3][6] = 16'b10100_000000_11111;
        onion_boiled[3][7] = 16'b10100_000000_11111;
        onion_boiled[3][8] = 16'b10100_000000_11111;
        onion_boiled[3][9] = 16'b10100_000000_11111;
        onion_boiled[3][10] = 16'b10100_000000_11111;
        onion_boiled[3][11] = 16'b11001_100101_11111;
        onion_boiled[3][12] = 16'b10100_000000_11111;
        onion_boiled[3][13] = 16'b00000_000000_00000;
        onion_boiled[3][14] = 16'b00000_000110_11111;
        onion_boiled[4][0] = 16'b00000_000110_11111;
        onion_boiled[4][1] = 16'b10100_000000_11111;
        onion_boiled[4][2] = 16'b11001_100101_11111;
        onion_boiled[4][3] = 16'b10100_000000_11111;
        onion_boiled[4][4] = 16'b10100_000000_11111;
        onion_boiled[4][5] = 16'b11001_100101_11111;
        onion_boiled[4][6] = 16'b11001_100101_11111;
        onion_boiled[4][7] = 16'b11001_100101_11111;
        onion_boiled[4][8] = 16'b11001_100101_11111;
        onion_boiled[4][9] = 16'b11001_100101_11111;
        onion_boiled[4][10] = 16'b10100_000000_11111;
        onion_boiled[4][11] = 16'b10100_000000_11111;
        onion_boiled[4][12] = 16'b11001_100101_11111;
        onion_boiled[4][13] = 16'b10100_000000_11111;
        onion_boiled[4][14] = 16'b00000_000110_11111;
        onion_boiled[5][0] = 16'b00000_000110_11111;
        onion_boiled[5][1] = 16'b10100_000000_11111;
        onion_boiled[5][2] = 16'b11001_100101_11111;
        onion_boiled[5][3] = 16'b10100_000000_11111;
        onion_boiled[5][4] = 16'b11001_100101_11111;
        onion_boiled[5][5] = 16'b10100_000000_11111;
        onion_boiled[5][6] = 16'b10100_000000_11111;
        onion_boiled[5][7] = 16'b10100_000000_11111;
        onion_boiled[5][8] = 16'b10100_000000_11111;
        onion_boiled[5][9] = 16'b10100_000000_11111;
        onion_boiled[5][10] = 16'b11001_100101_11111;
        onion_boiled[5][11] = 16'b10100_000000_11111;
        onion_boiled[5][12] = 16'b11001_100101_11111;
        onion_boiled[5][13] = 16'b10100_000000_11111;
        onion_boiled[5][14] = 16'b00000_000110_11111;
        onion_boiled[6][0] = 16'b00000_000110_11111;
        onion_boiled[6][1] = 16'b10100_000000_11111;
        onion_boiled[6][2] = 16'b11001_100101_11111;
        onion_boiled[6][3] = 16'b10100_000000_11111;
        onion_boiled[6][4] = 16'b11001_100101_11111;
        onion_boiled[6][5] = 16'b10100_000000_11111;
        onion_boiled[6][6] = 16'b10100_000000_11111;
        onion_boiled[6][7] = 16'b11001_100101_11111;
        onion_boiled[6][8] = 16'b10100_000000_11111;
        onion_boiled[6][9] = 16'b10100_000000_11111;
        onion_boiled[6][10] = 16'b11001_100101_11111;
        onion_boiled[6][11] = 16'b10100_000000_11111;
        onion_boiled[6][12] = 16'b11001_100101_11111;
        onion_boiled[6][13] = 16'b10100_000000_11111;
        onion_boiled[6][14] = 16'b00000_000110_11111;
        onion_boiled[7][0] = 16'b00000_000110_11111;
        onion_boiled[7][1] = 16'b00000_000000_00000;
        onion_boiled[7][2] = 16'b11001_100101_11111;
        onion_boiled[7][3] = 16'b10100_000000_11111;
        onion_boiled[7][4] = 16'b10100_000000_11111;
        onion_boiled[7][5] = 16'b11001_100101_11111;
        onion_boiled[7][6] = 16'b10100_000000_11111;
        onion_boiled[7][7] = 16'b10100_000000_11111;
        onion_boiled[7][8] = 16'b11001_100101_11111;
        onion_boiled[7][9] = 16'b10100_000000_11111;
        onion_boiled[7][10] = 16'b11001_100101_11111;
        onion_boiled[7][11] = 16'b10100_000000_11111;
        onion_boiled[7][12] = 16'b11001_100101_11111;
        onion_boiled[7][13] = 16'b10100_000000_11111;
        onion_boiled[7][14] = 16'b00000_000110_11111;
        onion_boiled[8][0] = 16'b00000_000110_11111;
        onion_boiled[8][1] = 16'b00000_000000_00000;
        onion_boiled[8][2] = 16'b10100_000000_11111;
        onion_boiled[8][3] = 16'b11001_100101_11111;
        onion_boiled[8][4] = 16'b10100_000000_11111;
        onion_boiled[8][5] = 16'b10100_000000_11111;
        onion_boiled[8][6] = 16'b11001_100101_11111;
        onion_boiled[8][7] = 16'b10100_000000_11111;
        onion_boiled[8][8] = 16'b10100_000000_11111;
        onion_boiled[8][9] = 16'b11001_100101_11111;
        onion_boiled[8][10] = 16'b10100_000000_11111;
        onion_boiled[8][11] = 16'b10100_000000_11111;
        onion_boiled[8][12] = 16'b11001_100101_11111;
        onion_boiled[8][13] = 16'b10100_000000_11111;
        onion_boiled[8][14] = 16'b00000_000110_11111;
        onion_boiled[9][0] = 16'b00000_000110_11111;
        onion_boiled[9][1] = 16'b00000_000000_00000;
        onion_boiled[9][2] = 16'b00000_000000_00000;
        onion_boiled[9][3] = 16'b10100_000000_11111;
        onion_boiled[9][4] = 16'b11001_100101_11111;
        onion_boiled[9][5] = 16'b10100_000000_11111;
        onion_boiled[9][6] = 16'b10100_000000_11111;
        onion_boiled[9][7] = 16'b11001_100101_11111;
        onion_boiled[9][8] = 16'b11001_100101_11111;
        onion_boiled[9][9] = 16'b10100_000000_11111;
        onion_boiled[9][10] = 16'b10100_000000_11111;
        onion_boiled[9][11] = 16'b11001_100101_11111;
        onion_boiled[9][12] = 16'b10100_000000_11111;
        onion_boiled[9][13] = 16'b00000_000000_00000;
        onion_boiled[9][14] = 16'b00000_000110_11111;
        onion_boiled[10][0] = 16'b00000_000110_11111;
        onion_boiled[10][1] = 16'b00000_000000_00000;
        onion_boiled[10][2] = 16'b00000_000000_00000;
        onion_boiled[10][3] = 16'b00000_000000_00000;
        onion_boiled[10][4] = 16'b10100_000000_11111;
        onion_boiled[10][5] = 16'b11001_100101_11111;
        onion_boiled[10][6] = 16'b10100_000000_11111;
        onion_boiled[10][7] = 16'b10100_000000_11111;
        onion_boiled[10][8] = 16'b10100_000000_11111;
        onion_boiled[10][9] = 16'b10100_000000_11111;
        onion_boiled[10][10] = 16'b11001_100101_11111;
        onion_boiled[10][11] = 16'b10100_000000_11111;
        onion_boiled[10][12] = 16'b00000_000000_00000;
        onion_boiled[10][13] = 16'b00000_000000_00000;
        onion_boiled[10][14] = 16'b00000_000110_11111;
        onion_boiled[11][0] = 16'b00000_000110_11111;
        onion_boiled[11][1] = 16'b00000_000000_00000;
        onion_boiled[11][2] = 16'b00000_000000_00000;
        onion_boiled[11][3] = 16'b00000_000000_00000;
        onion_boiled[11][4] = 16'b00000_000000_00000;
        onion_boiled[11][5] = 16'b10100_000000_11111;
        onion_boiled[11][6] = 16'b11001_100101_11111;
        onion_boiled[11][7] = 16'b10100_000000_11111;
        onion_boiled[11][8] = 16'b10100_000000_11111;
        onion_boiled[11][9] = 16'b11001_100101_11111;
        onion_boiled[11][10] = 16'b10100_000000_11111;
        onion_boiled[11][11] = 16'b00000_000000_00000;
        onion_boiled[11][12] = 16'b00000_000000_00000;
        onion_boiled[11][13] = 16'b00000_000000_00000;
        onion_boiled[11][14] = 16'b00000_000110_11111;
        onion_boiled[12][0] = 16'b00000_000110_11111;
        onion_boiled[12][1] = 16'b00000_000000_00000;
        onion_boiled[12][2] = 16'b00000_000000_00000;
        onion_boiled[12][3] = 16'b00000_000000_00000;
        onion_boiled[12][4] = 16'b00000_000000_00000;
        onion_boiled[12][5] = 16'b00000_000000_00000;
        onion_boiled[12][6] = 16'b10100_000000_11111;
        onion_boiled[12][7] = 16'b11001_100101_11111;
        onion_boiled[12][8] = 16'b11001_100101_11111;
        onion_boiled[12][9] = 16'b10100_000000_11111;
        onion_boiled[12][10] = 16'b00000_000000_00000;
        onion_boiled[12][11] = 16'b00000_000000_00000;
        onion_boiled[12][12] = 16'b00000_000000_00000;
        onion_boiled[12][13] = 16'b00000_000000_00000;
        onion_boiled[12][14] = 16'b00000_000110_11111;
        onion_boiled[13][0] = 16'b00000_000110_11111;
        onion_boiled[13][1] = 16'b00000_000000_00000;
        onion_boiled[13][2] = 16'b00000_000000_00000;
        onion_boiled[13][3] = 16'b00000_000000_00000;
        onion_boiled[13][4] = 16'b00000_000000_00000;
        onion_boiled[13][5] = 16'b00000_000000_00000;
        onion_boiled[13][6] = 16'b00000_000000_00000;
        onion_boiled[13][7] = 16'b10100_000000_11111;
        onion_boiled[13][8] = 16'b00000_000000_00000;
        onion_boiled[13][9] = 16'b00000_000000_00000;
        onion_boiled[13][10] = 16'b00000_000000_00000;
        onion_boiled[13][11] = 16'b00000_000000_00000;
        onion_boiled[13][12] = 16'b00000_000000_00000;
        onion_boiled[13][13] = 16'b00000_000000_00000;
        onion_boiled[13][14] = 16'b00000_000110_11111;
        onion_boiled[14][0] = 16'b00000_000110_11111;
        onion_boiled[14][1] = 16'b00000_000110_11111;
        onion_boiled[14][2] = 16'b00000_000110_11111;
        onion_boiled[14][3] = 16'b00000_000110_11111;
        onion_boiled[14][4] = 16'b00000_000110_11111;
        onion_boiled[14][5] = 16'b00000_000110_11111;
        onion_boiled[14][6] = 16'b00000_000110_11111;
        onion_boiled[14][7] = 16'b00000_000110_11111;
        onion_boiled[14][8] = 16'b00000_000110_11111;
        onion_boiled[14][9] = 16'b00000_000110_11111;
        onion_boiled[14][10] = 16'b00000_000110_11111;
        onion_boiled[14][11] = 16'b00000_000110_11111;
        onion_boiled[14][12] = 16'b00000_000110_11111;
        onion_boiled[14][13] = 16'b00000_000110_11111;
        onion_boiled[14][14] = 16'b00000_000110_11111;


        onion_chopped[0][0] = 16'b00000_111111_00001;
        onion_chopped[0][1] = 16'b00000_111111_00001;
        onion_chopped[0][2] = 16'b00000_111111_00001;
        onion_chopped[0][3] = 16'b00000_111111_00001;
        onion_chopped[0][4] = 16'b00000_111111_00001;
        onion_chopped[0][5] = 16'b00000_111111_00001;
        onion_chopped[0][6] = 16'b00000_111111_00001;
        onion_chopped[0][7] = 16'b00000_111111_00001;
        onion_chopped[0][8] = 16'b00000_111111_00001;
        onion_chopped[0][9] = 16'b00000_111111_00001;
        onion_chopped[0][10] = 16'b00000_111111_00001;
        onion_chopped[0][11] = 16'b00000_111111_00001;
        onion_chopped[0][12] = 16'b00000_111111_00001;
        onion_chopped[0][13] = 16'b00000_111111_00001;
        onion_chopped[0][14] = 16'b00000_111111_00001;
        onion_chopped[1][0] = 16'b00000_111111_00001;
        onion_chopped[1][1] = 16'b00000_000000_00000;
        onion_chopped[1][2] = 16'b00000_000000_00000;
        onion_chopped[1][3] = 16'b10100_000000_11111;
        onion_chopped[1][4] = 16'b10100_000000_11111;
        onion_chopped[1][5] = 16'b10100_000000_11111;
        onion_chopped[1][6] = 16'b10100_000000_11111;
        onion_chopped[1][7] = 16'b10100_000000_11111;
        onion_chopped[1][8] = 16'b10100_000000_11111;
        onion_chopped[1][9] = 16'b10100_000000_11111;
        onion_chopped[1][10] = 16'b10100_000000_11111;
        onion_chopped[1][11] = 16'b00000_000000_00000;
        onion_chopped[1][12] = 16'b00000_000000_00000;
        onion_chopped[1][13] = 16'b00000_000000_00000;
        onion_chopped[1][14] = 16'b00000_111111_00001;
        onion_chopped[2][0] = 16'b00000_111111_00001;
        onion_chopped[2][1] = 16'b00000_000000_00000;
        onion_chopped[2][2] = 16'b10100_000000_11111;
        onion_chopped[2][3] = 16'b10100_000000_11111;
        onion_chopped[2][4] = 16'b11001_100101_11111;
        onion_chopped[2][5] = 16'b11001_100101_11111;
        onion_chopped[2][6] = 16'b11001_100101_11111;
        onion_chopped[2][7] = 16'b11001_100101_11111;
        onion_chopped[2][8] = 16'b11001_100101_11111;
        onion_chopped[2][9] = 16'b11001_100101_11111;
        onion_chopped[2][10] = 16'b11001_100101_11111;
        onion_chopped[2][11] = 16'b11001_100101_11111;
        onion_chopped[2][12] = 16'b10100_000000_11111;
        onion_chopped[2][13] = 16'b00000_000000_00000;
        onion_chopped[2][14] = 16'b00000_111111_00001;
        onion_chopped[3][0] = 16'b00000_111111_00001;
        onion_chopped[3][1] = 16'b10100_000000_11111;
        onion_chopped[3][2] = 16'b10100_000000_11111;
        onion_chopped[3][3] = 16'b11001_100101_11111;
        onion_chopped[3][4] = 16'b10100_000000_11111;
        onion_chopped[3][5] = 16'b10100_000000_11111;
        onion_chopped[3][6] = 16'b10100_000000_11111;
        onion_chopped[3][7] = 16'b10100_000000_11111;
        onion_chopped[3][8] = 16'b10100_000000_11111;
        onion_chopped[3][9] = 16'b10100_000000_11111;
        onion_chopped[3][10] = 16'b10100_000000_11111;
        onion_chopped[3][11] = 16'b11001_100101_11111;
        onion_chopped[3][12] = 16'b10100_000000_11111;
        onion_chopped[3][13] = 16'b00000_000000_00000;
        onion_chopped[3][14] = 16'b00000_111111_00001;
        onion_chopped[4][0] = 16'b00000_111111_00001;
        onion_chopped[4][1] = 16'b10100_000000_11111;
        onion_chopped[4][2] = 16'b11001_100101_11111;
        onion_chopped[4][3] = 16'b10100_000000_11111;
        onion_chopped[4][4] = 16'b10100_000000_11111;
        onion_chopped[4][5] = 16'b11001_100101_11111;
        onion_chopped[4][6] = 16'b11001_100101_11111;
        onion_chopped[4][7] = 16'b11001_100101_11111;
        onion_chopped[4][8] = 16'b11001_100101_11111;
        onion_chopped[4][9] = 16'b11001_100101_11111;
        onion_chopped[4][10] = 16'b10100_000000_11111;
        onion_chopped[4][11] = 16'b10100_000000_11111;
        onion_chopped[4][12] = 16'b11001_100101_11111;
        onion_chopped[4][13] = 16'b10100_000000_11111;
        onion_chopped[4][14] = 16'b00000_111111_00001;
        onion_chopped[5][0] = 16'b00000_111111_00001;
        onion_chopped[5][1] = 16'b10100_000000_11111;
        onion_chopped[5][2] = 16'b11001_100101_11111;
        onion_chopped[5][3] = 16'b10100_000000_11111;
        onion_chopped[5][4] = 16'b11001_100101_11111;
        onion_chopped[5][5] = 16'b10100_000000_11111;
        onion_chopped[5][6] = 16'b10100_000000_11111;
        onion_chopped[5][7] = 16'b10100_000000_11111;
        onion_chopped[5][8] = 16'b10100_000000_11111;
        onion_chopped[5][9] = 16'b10100_000000_11111;
        onion_chopped[5][10] = 16'b11001_100101_11111;
        onion_chopped[5][11] = 16'b10100_000000_11111;
        onion_chopped[5][12] = 16'b11001_100101_11111;
        onion_chopped[5][13] = 16'b10100_000000_11111;
        onion_chopped[5][14] = 16'b00000_111111_00001;
        onion_chopped[6][0] = 16'b00000_111111_00001;
        onion_chopped[6][1] = 16'b10100_000000_11111;
        onion_chopped[6][2] = 16'b11001_100101_11111;
        onion_chopped[6][3] = 16'b10100_000000_11111;
        onion_chopped[6][4] = 16'b11001_100101_11111;
        onion_chopped[6][5] = 16'b10100_000000_11111;
        onion_chopped[6][6] = 16'b10100_000000_11111;
        onion_chopped[6][7] = 16'b11001_100101_11111;
        onion_chopped[6][8] = 16'b10100_000000_11111;
        onion_chopped[6][9] = 16'b10100_000000_11111;
        onion_chopped[6][10] = 16'b11001_100101_11111;
        onion_chopped[6][11] = 16'b10100_000000_11111;
        onion_chopped[6][12] = 16'b11001_100101_11111;
        onion_chopped[6][13] = 16'b10100_000000_11111;
        onion_chopped[6][14] = 16'b00000_111111_00001;
        onion_chopped[7][0] = 16'b00000_111111_00001;
        onion_chopped[7][1] = 16'b00000_000000_00000;
        onion_chopped[7][2] = 16'b11001_100101_11111;
        onion_chopped[7][3] = 16'b10100_000000_11111;
        onion_chopped[7][4] = 16'b10100_000000_11111;
        onion_chopped[7][5] = 16'b11001_100101_11111;
        onion_chopped[7][6] = 16'b10100_000000_11111;
        onion_chopped[7][7] = 16'b10100_000000_11111;
        onion_chopped[7][8] = 16'b11001_100101_11111;
        onion_chopped[7][9] = 16'b10100_000000_11111;
        onion_chopped[7][10] = 16'b11001_100101_11111;
        onion_chopped[7][11] = 16'b10100_000000_11111;
        onion_chopped[7][12] = 16'b11001_100101_11111;
        onion_chopped[7][13] = 16'b10100_000000_11111;
        onion_chopped[7][14] = 16'b00000_111111_00001;
        onion_chopped[8][0] = 16'b00000_111111_00001;
        onion_chopped[8][1] = 16'b00000_000000_00000;
        onion_chopped[8][2] = 16'b10100_000000_11111;
        onion_chopped[8][3] = 16'b11001_100101_11111;
        onion_chopped[8][4] = 16'b10100_000000_11111;
        onion_chopped[8][5] = 16'b10100_000000_11111;
        onion_chopped[8][6] = 16'b11001_100101_11111;
        onion_chopped[8][7] = 16'b10100_000000_11111;
        onion_chopped[8][8] = 16'b10100_000000_11111;
        onion_chopped[8][9] = 16'b11001_100101_11111;
        onion_chopped[8][10] = 16'b10100_000000_11111;
        onion_chopped[8][11] = 16'b10100_000000_11111;
        onion_chopped[8][12] = 16'b11001_100101_11111;
        onion_chopped[8][13] = 16'b10100_000000_11111;
        onion_chopped[8][14] = 16'b00000_111111_00001;
        onion_chopped[9][0] = 16'b00000_111111_00001;
        onion_chopped[9][1] = 16'b00000_000000_00000;
        onion_chopped[9][2] = 16'b00000_000000_00000;
        onion_chopped[9][3] = 16'b10100_000000_11111;
        onion_chopped[9][4] = 16'b11001_100101_11111;
        onion_chopped[9][5] = 16'b10100_000000_11111;
        onion_chopped[9][6] = 16'b10100_000000_11111;
        onion_chopped[9][7] = 16'b11001_100101_11111;
        onion_chopped[9][8] = 16'b11001_100101_11111;
        onion_chopped[9][9] = 16'b10100_000000_11111;
        onion_chopped[9][10] = 16'b10100_000000_11111;
        onion_chopped[9][11] = 16'b11001_100101_11111;
        onion_chopped[9][12] = 16'b10100_000000_11111;
        onion_chopped[9][13] = 16'b00000_000000_00000;
        onion_chopped[9][14] = 16'b00000_111111_00001;
        onion_chopped[10][0] = 16'b00000_111111_00001;
        onion_chopped[10][1] = 16'b00000_000000_00000;
        onion_chopped[10][2] = 16'b00000_000000_00000;
        onion_chopped[10][3] = 16'b00000_000000_00000;
        onion_chopped[10][4] = 16'b10100_000000_11111;
        onion_chopped[10][5] = 16'b11001_100101_11111;
        onion_chopped[10][6] = 16'b10100_000000_11111;
        onion_chopped[10][7] = 16'b10100_000000_11111;
        onion_chopped[10][8] = 16'b10100_000000_11111;
        onion_chopped[10][9] = 16'b10100_000000_11111;
        onion_chopped[10][10] = 16'b11001_100101_11111;
        onion_chopped[10][11] = 16'b10100_000000_11111;
        onion_chopped[10][12] = 16'b00000_000000_00000;
        onion_chopped[10][13] = 16'b00000_000000_00000;
        onion_chopped[10][14] = 16'b00000_111111_00001;
        onion_chopped[11][0] = 16'b00000_111111_00001;
        onion_chopped[11][1] = 16'b00000_000000_00000;
        onion_chopped[11][2] = 16'b00000_000000_00000;
        onion_chopped[11][3] = 16'b00000_000000_00000;
        onion_chopped[11][4] = 16'b00000_000000_00000;
        onion_chopped[11][5] = 16'b10100_000000_11111;
        onion_chopped[11][6] = 16'b11001_100101_11111;
        onion_chopped[11][7] = 16'b10100_000000_11111;
        onion_chopped[11][8] = 16'b10100_000000_11111;
        onion_chopped[11][9] = 16'b11001_100101_11111;
        onion_chopped[11][10] = 16'b10100_000000_11111;
        onion_chopped[11][11] = 16'b00000_000000_00000;
        onion_chopped[11][12] = 16'b00000_000000_00000;
        onion_chopped[11][13] = 16'b00000_000000_00000;
        onion_chopped[11][14] = 16'b00000_111111_00001;
        onion_chopped[12][0] = 16'b00000_111111_00001;
        onion_chopped[12][1] = 16'b00000_000000_00000;
        onion_chopped[12][2] = 16'b00000_000000_00000;
        onion_chopped[12][3] = 16'b00000_000000_00000;
        onion_chopped[12][4] = 16'b00000_000000_00000;
        onion_chopped[12][5] = 16'b00000_000000_00000;
        onion_chopped[12][6] = 16'b10100_000000_11111;
        onion_chopped[12][7] = 16'b11001_100101_11111;
        onion_chopped[12][8] = 16'b11001_100101_11111;
        onion_chopped[12][9] = 16'b10100_000000_11111;
        onion_chopped[12][10] = 16'b00000_000000_00000;
        onion_chopped[12][11] = 16'b00000_000000_00000;
        onion_chopped[12][12] = 16'b00000_000000_00000;
        onion_chopped[12][13] = 16'b00000_000000_00000;
        onion_chopped[12][14] = 16'b00000_111111_00001;
        onion_chopped[13][0] = 16'b00000_111111_00001;
        onion_chopped[13][1] = 16'b00000_000000_00000;
        onion_chopped[13][2] = 16'b00000_000000_00000;
        onion_chopped[13][3] = 16'b00000_000000_00000;
        onion_chopped[13][4] = 16'b00000_000000_00000;
        onion_chopped[13][5] = 16'b00000_000000_00000;
        onion_chopped[13][6] = 16'b00000_000000_00000;
        onion_chopped[13][7] = 16'b10100_000000_11111;
        onion_chopped[13][8] = 16'b00000_000000_00000;
        onion_chopped[13][9] = 16'b00000_000000_00000;
        onion_chopped[13][10] = 16'b00000_000000_00000;
        onion_chopped[13][11] = 16'b00000_000000_00000;
        onion_chopped[13][12] = 16'b00000_000000_00000;
        onion_chopped[13][13] = 16'b00000_000000_00000;
        onion_chopped[13][14] = 16'b00000_111111_00001;
        onion_chopped[14][0] = 16'b00000_111111_00001;
        onion_chopped[14][1] = 16'b00000_111111_00001;
        onion_chopped[14][2] = 16'b00000_111111_00001;
        onion_chopped[14][3] = 16'b00000_111111_00001;
        onion_chopped[14][4] = 16'b00000_111111_00001;
        onion_chopped[14][5] = 16'b00000_111111_00001;
        onion_chopped[14][6] = 16'b00000_111111_00001;
        onion_chopped[14][7] = 16'b00000_111111_00001;
        onion_chopped[14][8] = 16'b00000_111111_00001;
        onion_chopped[14][9] = 16'b00000_111111_00001;
        onion_chopped[14][10] = 16'b00000_111111_00001;
        onion_chopped[14][11] = 16'b00000_111111_00001;
        onion_chopped[14][12] = 16'b00000_111111_00001;
        onion_chopped[14][13] = 16'b00000_111111_00001;
        onion_chopped[14][14] = 16'b00000_111111_00001;


        onion_raw[0][0] = 16'b11001_100101_11111;
        onion_raw[0][1] = 16'b11001_100101_11111;
        onion_raw[0][2] = 16'b11001_100101_11111;
        onion_raw[0][3] = 16'b11001_100101_11111;
        onion_raw[0][4] = 16'b11001_100101_11111;
        onion_raw[0][5] = 16'b11001_100101_11111;
        onion_raw[0][6] = 16'b11001_100101_11111;
        onion_raw[0][7] = 16'b11001_100101_11111;
        onion_raw[0][8] = 16'b11001_100101_11111;
        onion_raw[0][9] = 16'b11001_100101_11111;
        onion_raw[0][10] = 16'b11001_100101_11111;
        onion_raw[0][11] = 16'b11001_100101_11111;
        onion_raw[0][12] = 16'b11001_100101_11111;
        onion_raw[0][13] = 16'b11001_100101_11111;
        onion_raw[0][14] = 16'b11001_100101_11111;
        onion_raw[1][0] = 16'b11001_100101_11111;
        onion_raw[1][1] = 16'b00000_000000_00000;
        onion_raw[1][2] = 16'b00000_000000_00000;
        onion_raw[1][3] = 16'b10100_000000_11111;
        onion_raw[1][4] = 16'b10100_000000_11111;
        onion_raw[1][5] = 16'b10100_000000_11111;
        onion_raw[1][6] = 16'b10100_000000_11111;
        onion_raw[1][7] = 16'b10100_000000_11111;
        onion_raw[1][8] = 16'b10100_000000_11111;
        onion_raw[1][9] = 16'b10100_000000_11111;
        onion_raw[1][10] = 16'b10100_000000_11111;
        onion_raw[1][11] = 16'b00000_000000_00000;
        onion_raw[1][12] = 16'b00000_000000_00000;
        onion_raw[1][13] = 16'b00000_000000_00000;
        onion_raw[1][14] = 16'b11001_100101_11111;
        onion_raw[2][0] = 16'b11001_100101_11111;
        onion_raw[2][1] = 16'b00000_000000_00000;
        onion_raw[2][2] = 16'b10100_000000_11111;
        onion_raw[2][3] = 16'b10100_000000_11111;
        onion_raw[2][4] = 16'b11001_100101_11111;
        onion_raw[2][5] = 16'b11001_100101_11111;
        onion_raw[2][6] = 16'b11001_100101_11111;
        onion_raw[2][7] = 16'b11001_100101_11111;
        onion_raw[2][8] = 16'b11001_100101_11111;
        onion_raw[2][9] = 16'b11001_100101_11111;
        onion_raw[2][10] = 16'b11001_100101_11111;
        onion_raw[2][11] = 16'b11001_100101_11111;
        onion_raw[2][12] = 16'b10100_000000_11111;
        onion_raw[2][13] = 16'b00000_000000_00000;
        onion_raw[2][14] = 16'b11001_100101_11111;
        onion_raw[3][0] = 16'b11001_100101_11111;
        onion_raw[3][1] = 16'b10100_000000_11111;
        onion_raw[3][2] = 16'b10100_000000_11111;
        onion_raw[3][3] = 16'b11001_100101_11111;
        onion_raw[3][4] = 16'b10100_000000_11111;
        onion_raw[3][5] = 16'b10100_000000_11111;
        onion_raw[3][6] = 16'b10100_000000_11111;
        onion_raw[3][7] = 16'b10100_000000_11111;
        onion_raw[3][8] = 16'b10100_000000_11111;
        onion_raw[3][9] = 16'b10100_000000_11111;
        onion_raw[3][10] = 16'b10100_000000_11111;
        onion_raw[3][11] = 16'b11001_100101_11111;
        onion_raw[3][12] = 16'b10100_000000_11111;
        onion_raw[3][13] = 16'b00000_000000_00000;
        onion_raw[3][14] = 16'b11001_100101_11111;
        onion_raw[4][0] = 16'b11001_100101_11111;
        onion_raw[4][1] = 16'b10100_000000_11111;
        onion_raw[4][2] = 16'b11001_100101_11111;
        onion_raw[4][3] = 16'b10100_000000_11111;
        onion_raw[4][4] = 16'b10100_000000_11111;
        onion_raw[4][5] = 16'b11001_100101_11111;
        onion_raw[4][6] = 16'b11001_100101_11111;
        onion_raw[4][7] = 16'b11001_100101_11111;
        onion_raw[4][8] = 16'b11001_100101_11111;
        onion_raw[4][9] = 16'b11001_100101_11111;
        onion_raw[4][10] = 16'b10100_000000_11111;
        onion_raw[4][11] = 16'b10100_000000_11111;
        onion_raw[4][12] = 16'b11001_100101_11111;
        onion_raw[4][13] = 16'b10100_000000_11111;
        onion_raw[4][14] = 16'b11001_100101_11111;
        onion_raw[5][0] = 16'b11001_100101_11111;
        onion_raw[5][1] = 16'b10100_000000_11111;
        onion_raw[5][2] = 16'b11001_100101_11111;
        onion_raw[5][3] = 16'b10100_000000_11111;
        onion_raw[5][4] = 16'b11001_100101_11111;
        onion_raw[5][5] = 16'b10100_000000_11111;
        onion_raw[5][6] = 16'b10100_000000_11111;
        onion_raw[5][7] = 16'b10100_000000_11111;
        onion_raw[5][8] = 16'b10100_000000_11111;
        onion_raw[5][9] = 16'b10100_000000_11111;
        onion_raw[5][10] = 16'b11001_100101_11111;
        onion_raw[5][11] = 16'b10100_000000_11111;
        onion_raw[5][12] = 16'b11001_100101_11111;
        onion_raw[5][13] = 16'b10100_000000_11111;
        onion_raw[5][14] = 16'b11001_100101_11111;
        onion_raw[6][0] = 16'b11001_100101_11111;
        onion_raw[6][1] = 16'b10100_000000_11111;
        onion_raw[6][2] = 16'b11001_100101_11111;
        onion_raw[6][3] = 16'b10100_000000_11111;
        onion_raw[6][4] = 16'b11001_100101_11111;
        onion_raw[6][5] = 16'b10100_000000_11111;
        onion_raw[6][6] = 16'b10100_000000_11111;
        onion_raw[6][7] = 16'b11001_100101_11111;
        onion_raw[6][8] = 16'b10100_000000_11111;
        onion_raw[6][9] = 16'b10100_000000_11111;
        onion_raw[6][10] = 16'b11001_100101_11111;
        onion_raw[6][11] = 16'b10100_000000_11111;
        onion_raw[6][12] = 16'b11001_100101_11111;
        onion_raw[6][13] = 16'b10100_000000_11111;
        onion_raw[6][14] = 16'b11001_100101_11111;
        onion_raw[7][0] = 16'b11001_100101_11111;
        onion_raw[7][1] = 16'b00000_000000_00000;
        onion_raw[7][2] = 16'b11001_100101_11111;
        onion_raw[7][3] = 16'b10100_000000_11111;
        onion_raw[7][4] = 16'b10100_000000_11111;
        onion_raw[7][5] = 16'b11001_100101_11111;
        onion_raw[7][6] = 16'b10100_000000_11111;
        onion_raw[7][7] = 16'b10100_000000_11111;
        onion_raw[7][8] = 16'b11001_100101_11111;
        onion_raw[7][9] = 16'b10100_000000_11111;
        onion_raw[7][10] = 16'b11001_100101_11111;
        onion_raw[7][11] = 16'b10100_000000_11111;
        onion_raw[7][12] = 16'b11001_100101_11111;
        onion_raw[7][13] = 16'b10100_000000_11111;
        onion_raw[7][14] = 16'b11001_100101_11111;
        onion_raw[8][0] = 16'b11001_100101_11111;
        onion_raw[8][1] = 16'b00000_000000_00000;
        onion_raw[8][2] = 16'b10100_000000_11111;
        onion_raw[8][3] = 16'b11001_100101_11111;
        onion_raw[8][4] = 16'b10100_000000_11111;
        onion_raw[8][5] = 16'b10100_000000_11111;
        onion_raw[8][6] = 16'b11001_100101_11111;
        onion_raw[8][7] = 16'b10100_000000_11111;
        onion_raw[8][8] = 16'b10100_000000_11111;
        onion_raw[8][9] = 16'b11001_100101_11111;
        onion_raw[8][10] = 16'b10100_000000_11111;
        onion_raw[8][11] = 16'b10100_000000_11111;
        onion_raw[8][12] = 16'b11001_100101_11111;
        onion_raw[8][13] = 16'b10100_000000_11111;
        onion_raw[8][14] = 16'b11001_100101_11111;
        onion_raw[9][0] = 16'b11001_100101_11111;
        onion_raw[9][1] = 16'b00000_000000_00000;
        onion_raw[9][2] = 16'b00000_000000_00000;
        onion_raw[9][3] = 16'b10100_000000_11111;
        onion_raw[9][4] = 16'b11001_100101_11111;
        onion_raw[9][5] = 16'b10100_000000_11111;
        onion_raw[9][6] = 16'b10100_000000_11111;
        onion_raw[9][7] = 16'b11001_100101_11111;
        onion_raw[9][8] = 16'b11001_100101_11111;
        onion_raw[9][9] = 16'b10100_000000_11111;
        onion_raw[9][10] = 16'b10100_000000_11111;
        onion_raw[9][11] = 16'b11001_100101_11111;
        onion_raw[9][12] = 16'b10100_000000_11111;
        onion_raw[9][13] = 16'b00000_000000_00000;
        onion_raw[9][14] = 16'b11001_100101_11111;
        onion_raw[10][0] = 16'b11001_100101_11111;
        onion_raw[10][1] = 16'b00000_000000_00000;
        onion_raw[10][2] = 16'b00000_000000_00000;
        onion_raw[10][3] = 16'b00000_000000_00000;
        onion_raw[10][4] = 16'b10100_000000_11111;
        onion_raw[10][5] = 16'b11001_100101_11111;
        onion_raw[10][6] = 16'b10100_000000_11111;
        onion_raw[10][7] = 16'b10100_000000_11111;
        onion_raw[10][8] = 16'b10100_000000_11111;
        onion_raw[10][9] = 16'b10100_000000_11111;
        onion_raw[10][10] = 16'b11001_100101_11111;
        onion_raw[10][11] = 16'b10100_000000_11111;
        onion_raw[10][12] = 16'b00000_000000_00000;
        onion_raw[10][13] = 16'b00000_000000_00000;
        onion_raw[10][14] = 16'b11001_100101_11111;
        onion_raw[11][0] = 16'b11001_100101_11111;
        onion_raw[11][1] = 16'b00000_000000_00000;
        onion_raw[11][2] = 16'b00000_000000_00000;
        onion_raw[11][3] = 16'b00000_000000_00000;
        onion_raw[11][4] = 16'b00000_000000_00000;
        onion_raw[11][5] = 16'b10100_000000_11111;
        onion_raw[11][6] = 16'b11001_100101_11111;
        onion_raw[11][7] = 16'b10100_000000_11111;
        onion_raw[11][8] = 16'b10100_000000_11111;
        onion_raw[11][9] = 16'b11001_100101_11111;
        onion_raw[11][10] = 16'b10100_000000_11111;
        onion_raw[11][11] = 16'b00000_000000_00000;
        onion_raw[11][12] = 16'b00000_000000_00000;
        onion_raw[11][13] = 16'b00000_000000_00000;
        onion_raw[11][14] = 16'b11001_100101_11111;
        onion_raw[12][0] = 16'b11001_100101_11111;
        onion_raw[12][1] = 16'b00000_000000_00000;
        onion_raw[12][2] = 16'b00000_000000_00000;
        onion_raw[12][3] = 16'b00000_000000_00000;
        onion_raw[12][4] = 16'b00000_000000_00000;
        onion_raw[12][5] = 16'b00000_000000_00000;
        onion_raw[12][6] = 16'b10100_000000_11111;
        onion_raw[12][7] = 16'b11001_100101_11111;
        onion_raw[12][8] = 16'b11001_100101_11111;
        onion_raw[12][9] = 16'b10100_000000_11111;
        onion_raw[12][10] = 16'b00000_000000_00000;
        onion_raw[12][11] = 16'b00000_000000_00000;
        onion_raw[12][12] = 16'b00000_000000_00000;
        onion_raw[12][13] = 16'b00000_000000_00000;
        onion_raw[12][14] = 16'b11001_100101_11111;
        onion_raw[13][0] = 16'b11001_100101_11111;
        onion_raw[13][1] = 16'b00000_000000_00000;
        onion_raw[13][2] = 16'b00000_000000_00000;
        onion_raw[13][3] = 16'b00000_000000_00000;
        onion_raw[13][4] = 16'b00000_000000_00000;
        onion_raw[13][5] = 16'b00000_000000_00000;
        onion_raw[13][6] = 16'b00000_000000_00000;
        onion_raw[13][7] = 16'b10100_000000_11111;
        onion_raw[13][8] = 16'b00000_000000_00000;
        onion_raw[13][9] = 16'b00000_000000_00000;
        onion_raw[13][10] = 16'b00000_000000_00000;
        onion_raw[13][11] = 16'b00000_000000_00000;
        onion_raw[13][12] = 16'b00000_000000_00000;
        onion_raw[13][13] = 16'b00000_000000_00000;
        onion_raw[13][14] = 16'b11001_100101_11111;
        onion_raw[14][0] = 16'b11001_100101_11111;
        onion_raw[14][1] = 16'b11001_100101_11111;
        onion_raw[14][2] = 16'b11001_100101_11111;
        onion_raw[14][3] = 16'b11001_100101_11111;
        onion_raw[14][4] = 16'b11001_100101_11111;
        onion_raw[14][5] = 16'b11001_100101_11111;
        onion_raw[14][6] = 16'b11001_100101_11111;
        onion_raw[14][7] = 16'b11001_100101_11111;
        onion_raw[14][8] = 16'b11001_100101_11111;
        onion_raw[14][9] = 16'b11001_100101_11111;
        onion_raw[14][10] = 16'b11001_100101_11111;
        onion_raw[14][11] = 16'b11001_100101_11111;
        onion_raw[14][12] = 16'b11001_100101_11111;
        onion_raw[14][13] = 16'b11001_100101_11111;
        onion_raw[14][14] = 16'b11001_100101_11111;


        tomato_boiled_chopped[0][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][1] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][2] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][3] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][4] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][5] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][6] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][7] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][8] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][9] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][10] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][11] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][12] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][13] = 16'b10101_011000_00000;
        tomato_boiled_chopped[0][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[1][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[1][1] = 16'b00000_000000_00000;
        tomato_boiled_chopped[1][2] = 16'b00000_000000_00000;
        tomato_boiled_chopped[1][3] = 16'b00000_000000_00000;
        tomato_boiled_chopped[1][4] = 16'b00000_000000_00000;
        tomato_boiled_chopped[1][5] = 16'b00000_000000_00000;
        tomato_boiled_chopped[1][6] = 16'b00000_000000_00000;
        tomato_boiled_chopped[1][7] = 16'b00000_000000_00000;
        tomato_boiled_chopped[1][8] = 16'b00000_000000_00000;
        tomato_boiled_chopped[1][9] = 16'b00000_000000_00000;
        tomato_boiled_chopped[1][10] = 16'b00000_000000_00000;
        tomato_boiled_chopped[1][11] = 16'b00000_000000_00000;
        tomato_boiled_chopped[1][12] = 16'b00000_000000_00000;
        tomato_boiled_chopped[1][13] = 16'b00000_000000_00000;
        tomato_boiled_chopped[1][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[2][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[2][1] = 16'b00000_000000_00000;
        tomato_boiled_chopped[2][2] = 16'b00000_000000_00000;
        tomato_boiled_chopped[2][3] = 16'b00000_000000_00000;
        tomato_boiled_chopped[2][4] = 16'b00000_000000_00000;
        tomato_boiled_chopped[2][5] = 16'b10001_000000_00000;
        tomato_boiled_chopped[2][6] = 16'b10001_000000_00000;
        tomato_boiled_chopped[2][7] = 16'b10001_000000_00000;
        tomato_boiled_chopped[2][8] = 16'b10001_000000_00000;
        tomato_boiled_chopped[2][9] = 16'b10001_000000_00000;
        tomato_boiled_chopped[2][10] = 16'b00000_000000_00000;
        tomato_boiled_chopped[2][11] = 16'b00000_000000_00000;
        tomato_boiled_chopped[2][12] = 16'b00000_000000_00000;
        tomato_boiled_chopped[2][13] = 16'b00000_000000_00000;
        tomato_boiled_chopped[2][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[3][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[3][1] = 16'b00000_000000_00000;
        tomato_boiled_chopped[3][2] = 16'b00000_000000_00000;
        tomato_boiled_chopped[3][3] = 16'b10001_000000_00000;
        tomato_boiled_chopped[3][4] = 16'b10001_000000_00000;
        tomato_boiled_chopped[3][5] = 16'b10001_000000_00000;
        tomato_boiled_chopped[3][6] = 16'b11001_000000_00000;
        tomato_boiled_chopped[3][7] = 16'b11001_000000_00000;
        tomato_boiled_chopped[3][8] = 16'b11001_000000_00000;
        tomato_boiled_chopped[3][9] = 16'b10001_000000_00000;
        tomato_boiled_chopped[3][10] = 16'b10001_000000_00000;
        tomato_boiled_chopped[3][11] = 16'b10001_000000_00000;
        tomato_boiled_chopped[3][12] = 16'b00000_000000_00000;
        tomato_boiled_chopped[3][13] = 16'b00000_000000_00000;
        tomato_boiled_chopped[3][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[4][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[4][1] = 16'b00000_000000_00000;
        tomato_boiled_chopped[4][2] = 16'b10001_000000_00000;
        tomato_boiled_chopped[4][3] = 16'b11001_000000_00000;
        tomato_boiled_chopped[4][4] = 16'b11001_000000_00000;
        tomato_boiled_chopped[4][5] = 16'b11001_000000_00000;
        tomato_boiled_chopped[4][6] = 16'b11001_000000_00000;
        tomato_boiled_chopped[4][7] = 16'b11001_000000_00000;
        tomato_boiled_chopped[4][8] = 16'b11001_000000_00000;
        tomato_boiled_chopped[4][9] = 16'b11001_000000_00000;
        tomato_boiled_chopped[4][10] = 16'b11001_000000_00000;
        tomato_boiled_chopped[4][11] = 16'b11001_000000_00000;
        tomato_boiled_chopped[4][12] = 16'b10001_000000_00000;
        tomato_boiled_chopped[4][13] = 16'b00000_000000_00000;
        tomato_boiled_chopped[4][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[5][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[5][1] = 16'b00000_000000_00000;
        tomato_boiled_chopped[5][2] = 16'b11001_000000_00000;
        tomato_boiled_chopped[5][3] = 16'b11001_000000_00000;
        tomato_boiled_chopped[5][4] = 16'b11001_000000_00000;
        tomato_boiled_chopped[5][5] = 16'b11001_000000_00000;
        tomato_boiled_chopped[5][6] = 16'b11001_000000_00000;
        tomato_boiled_chopped[5][7] = 16'b11001_000000_00000;
        tomato_boiled_chopped[5][8] = 16'b11001_000000_00000;
        tomato_boiled_chopped[5][9] = 16'b11001_000000_00000;
        tomato_boiled_chopped[5][10] = 16'b11001_000000_00000;
        tomato_boiled_chopped[5][11] = 16'b11001_000000_00000;
        tomato_boiled_chopped[5][12] = 16'b11001_000000_00000;
        tomato_boiled_chopped[5][13] = 16'b00000_000000_00000;
        tomato_boiled_chopped[5][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[6][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[6][1] = 16'b00000_000000_00000;
        tomato_boiled_chopped[6][2] = 16'b11001_000000_00000;
        tomato_boiled_chopped[6][3] = 16'b11001_000000_00000;
        tomato_boiled_chopped[6][4] = 16'b11001_000000_00000;
        tomato_boiled_chopped[6][5] = 16'b11001_000000_00000;
        tomato_boiled_chopped[6][6] = 16'b11001_000000_00000;
        tomato_boiled_chopped[6][7] = 16'b11001_000000_00000;
        tomato_boiled_chopped[6][8] = 16'b11001_000000_00000;
        tomato_boiled_chopped[6][9] = 16'b11001_000000_00000;
        tomato_boiled_chopped[6][10] = 16'b11001_000000_00000;
        tomato_boiled_chopped[6][11] = 16'b11001_000000_00000;
        tomato_boiled_chopped[6][12] = 16'b11001_000000_00000;
        tomato_boiled_chopped[6][13] = 16'b00000_000000_00000;
        tomato_boiled_chopped[6][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[7][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[7][1] = 16'b00000_000000_00000;
        tomato_boiled_chopped[7][2] = 16'b11001_000000_00000;
        tomato_boiled_chopped[7][3] = 16'b11001_000000_00000;
        tomato_boiled_chopped[7][4] = 16'b11001_000000_00000;
        tomato_boiled_chopped[7][5] = 16'b11001_000000_00000;
        tomato_boiled_chopped[7][6] = 16'b11001_000000_00000;
        tomato_boiled_chopped[7][7] = 16'b11001_000000_00000;
        tomato_boiled_chopped[7][8] = 16'b11001_000000_00000;
        tomato_boiled_chopped[7][9] = 16'b11001_000000_00000;
        tomato_boiled_chopped[7][10] = 16'b11001_000000_00000;
        tomato_boiled_chopped[7][11] = 16'b11001_000000_00000;
        tomato_boiled_chopped[7][12] = 16'b11001_000000_00000;
        tomato_boiled_chopped[7][13] = 16'b00000_000000_00000;
        tomato_boiled_chopped[7][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[8][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[8][1] = 16'b00000_000000_00000;
        tomato_boiled_chopped[8][2] = 16'b11001_000000_00000;
        tomato_boiled_chopped[8][3] = 16'b00000_011100_00000;
        tomato_boiled_chopped[8][4] = 16'b11001_000000_00000;
        tomato_boiled_chopped[8][5] = 16'b11001_000000_00000;
        tomato_boiled_chopped[8][6] = 16'b11001_000000_00000;
        tomato_boiled_chopped[8][7] = 16'b11001_000000_00000;
        tomato_boiled_chopped[8][8] = 16'b11001_000000_00000;
        tomato_boiled_chopped[8][9] = 16'b11001_000000_00000;
        tomato_boiled_chopped[8][10] = 16'b11001_000000_00000;
        tomato_boiled_chopped[8][11] = 16'b00000_011100_00000;
        tomato_boiled_chopped[8][12] = 16'b11001_000000_00000;
        tomato_boiled_chopped[8][13] = 16'b00000_000000_00000;
        tomato_boiled_chopped[8][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[9][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[9][1] = 16'b00000_000000_00000;
        tomato_boiled_chopped[9][2] = 16'b11001_000000_00000;
        tomato_boiled_chopped[9][3] = 16'b00000_011100_00000;
        tomato_boiled_chopped[9][4] = 16'b00000_011100_00000;
        tomato_boiled_chopped[9][5] = 16'b00000_011100_00000;
        tomato_boiled_chopped[9][6] = 16'b11001_000000_00000;
        tomato_boiled_chopped[9][7] = 16'b11001_000000_00000;
        tomato_boiled_chopped[9][8] = 16'b11001_000000_00000;
        tomato_boiled_chopped[9][9] = 16'b00000_011100_00000;
        tomato_boiled_chopped[9][10] = 16'b00000_011100_00000;
        tomato_boiled_chopped[9][11] = 16'b00000_011100_00000;
        tomato_boiled_chopped[9][12] = 16'b11001_000000_00000;
        tomato_boiled_chopped[9][13] = 16'b00000_000000_00000;
        tomato_boiled_chopped[9][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[10][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[10][1] = 16'b00000_000000_00000;
        tomato_boiled_chopped[10][2] = 16'b00000_000000_00000;
        tomato_boiled_chopped[10][3] = 16'b11001_000000_00000;
        tomato_boiled_chopped[10][4] = 16'b00000_011100_00000;
        tomato_boiled_chopped[10][5] = 16'b00000_011100_00000;
        tomato_boiled_chopped[10][6] = 16'b00000_011100_00000;
        tomato_boiled_chopped[10][7] = 16'b11001_000000_00000;
        tomato_boiled_chopped[10][8] = 16'b00000_011100_00000;
        tomato_boiled_chopped[10][9] = 16'b00000_011100_00000;
        tomato_boiled_chopped[10][10] = 16'b00000_011100_00000;
        tomato_boiled_chopped[10][11] = 16'b11001_000000_00000;
        tomato_boiled_chopped[10][12] = 16'b00000_000000_00000;
        tomato_boiled_chopped[10][13] = 16'b00000_000000_00000;
        tomato_boiled_chopped[10][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[11][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[11][1] = 16'b00000_000000_00000;
        tomato_boiled_chopped[11][2] = 16'b00000_000000_00000;
        tomato_boiled_chopped[11][3] = 16'b00000_000000_00000;
        tomato_boiled_chopped[11][4] = 16'b11001_000000_00000;
        tomato_boiled_chopped[11][5] = 16'b11001_000000_00000;
        tomato_boiled_chopped[11][6] = 16'b00000_011100_00000;
        tomato_boiled_chopped[11][7] = 16'b00000_011100_00000;
        tomato_boiled_chopped[11][8] = 16'b00000_011100_00000;
        tomato_boiled_chopped[11][9] = 16'b11001_000000_00000;
        tomato_boiled_chopped[11][10] = 16'b11001_000000_00000;
        tomato_boiled_chopped[11][11] = 16'b00000_000000_00000;
        tomato_boiled_chopped[11][12] = 16'b00000_000000_00000;
        tomato_boiled_chopped[11][13] = 16'b00000_000000_00000;
        tomato_boiled_chopped[11][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[12][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[12][1] = 16'b00000_000000_00000;
        tomato_boiled_chopped[12][2] = 16'b00000_000000_00000;
        tomato_boiled_chopped[12][3] = 16'b00000_011100_00000;
        tomato_boiled_chopped[12][4] = 16'b00000_011100_00000;
        tomato_boiled_chopped[12][5] = 16'b00000_011100_00000;
        tomato_boiled_chopped[12][6] = 16'b00000_011100_00000;
        tomato_boiled_chopped[12][7] = 16'b11001_000000_00000;
        tomato_boiled_chopped[12][8] = 16'b00000_011100_00000;
        tomato_boiled_chopped[12][9] = 16'b00000_011100_00000;
        tomato_boiled_chopped[12][10] = 16'b00000_011100_00000;
        tomato_boiled_chopped[12][11] = 16'b00000_011100_00000;
        tomato_boiled_chopped[12][12] = 16'b00000_000000_00000;
        tomato_boiled_chopped[12][13] = 16'b00000_000000_00000;
        tomato_boiled_chopped[12][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[13][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[13][1] = 16'b00000_000000_00000;
        tomato_boiled_chopped[13][2] = 16'b00000_000000_00000;
        tomato_boiled_chopped[13][3] = 16'b00000_000000_00000;
        tomato_boiled_chopped[13][4] = 16'b00000_011100_00000;
        tomato_boiled_chopped[13][5] = 16'b00000_011100_00000;
        tomato_boiled_chopped[13][6] = 16'b00000_000000_00000;
        tomato_boiled_chopped[13][7] = 16'b00000_000000_00000;
        tomato_boiled_chopped[13][8] = 16'b00000_000000_00000;
        tomato_boiled_chopped[13][9] = 16'b00000_011100_00000;
        tomato_boiled_chopped[13][10] = 16'b00000_011100_00000;
        tomato_boiled_chopped[13][11] = 16'b00000_000000_00000;
        tomato_boiled_chopped[13][12] = 16'b00000_000000_00000;
        tomato_boiled_chopped[13][13] = 16'b00000_000000_00000;
        tomato_boiled_chopped[13][14] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][0] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][1] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][2] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][3] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][4] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][5] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][6] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][7] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][8] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][9] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][10] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][11] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][12] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][13] = 16'b10101_011000_00000;
        tomato_boiled_chopped[14][14] = 16'b10101_011000_00000;


        tomato_boiled[0][0] = 16'b00000_000110_11111;
        tomato_boiled[0][1] = 16'b00000_000110_11111;
        tomato_boiled[0][2] = 16'b00000_000110_11111;
        tomato_boiled[0][3] = 16'b00000_000110_11111;
        tomato_boiled[0][4] = 16'b00000_000110_11111;
        tomato_boiled[0][5] = 16'b00000_000110_11111;
        tomato_boiled[0][6] = 16'b00000_000110_11111;
        tomato_boiled[0][7] = 16'b00000_000110_11111;
        tomato_boiled[0][8] = 16'b00000_000110_11111;
        tomato_boiled[0][9] = 16'b00000_000110_11111;
        tomato_boiled[0][10] = 16'b00000_000110_11111;
        tomato_boiled[0][11] = 16'b00000_000110_11111;
        tomato_boiled[0][12] = 16'b00000_000110_11111;
        tomato_boiled[0][13] = 16'b00000_000110_11111;
        tomato_boiled[0][14] = 16'b00000_000110_11111;
        tomato_boiled[1][0] = 16'b00000_000110_11111;
        tomato_boiled[1][1] = 16'b00000_000000_00000;
        tomato_boiled[1][2] = 16'b00000_000000_00000;
        tomato_boiled[1][3] = 16'b00000_000000_00000;
        tomato_boiled[1][4] = 16'b00000_000000_00000;
        tomato_boiled[1][5] = 16'b00000_000000_00000;
        tomato_boiled[1][6] = 16'b00000_000000_00000;
        tomato_boiled[1][7] = 16'b00000_000000_00000;
        tomato_boiled[1][8] = 16'b00000_000000_00000;
        tomato_boiled[1][9] = 16'b00000_000000_00000;
        tomato_boiled[1][10] = 16'b00000_000000_00000;
        tomato_boiled[1][11] = 16'b00000_000000_00000;
        tomato_boiled[1][12] = 16'b00000_000000_00000;
        tomato_boiled[1][13] = 16'b00000_000000_00000;
        tomato_boiled[1][14] = 16'b00000_000110_11111;
        tomato_boiled[2][0] = 16'b00000_000110_11111;
        tomato_boiled[2][1] = 16'b00000_000000_00000;
        tomato_boiled[2][2] = 16'b00000_000000_00000;
        tomato_boiled[2][3] = 16'b00000_000000_00000;
        tomato_boiled[2][4] = 16'b00000_000000_00000;
        tomato_boiled[2][5] = 16'b10001_000000_00000;
        tomato_boiled[2][6] = 16'b10001_000000_00000;
        tomato_boiled[2][7] = 16'b10001_000000_00000;
        tomato_boiled[2][8] = 16'b10001_000000_00000;
        tomato_boiled[2][9] = 16'b10001_000000_00000;
        tomato_boiled[2][10] = 16'b00000_000000_00000;
        tomato_boiled[2][11] = 16'b00000_000000_00000;
        tomato_boiled[2][12] = 16'b00000_000000_00000;
        tomato_boiled[2][13] = 16'b00000_000000_00000;
        tomato_boiled[2][14] = 16'b00000_000110_11111;
        tomato_boiled[3][0] = 16'b00000_000110_11111;
        tomato_boiled[3][1] = 16'b00000_000000_00000;
        tomato_boiled[3][2] = 16'b00000_000000_00000;
        tomato_boiled[3][3] = 16'b10001_000000_00000;
        tomato_boiled[3][4] = 16'b10001_000000_00000;
        tomato_boiled[3][5] = 16'b10001_000000_00000;
        tomato_boiled[3][6] = 16'b11001_000000_00000;
        tomato_boiled[3][7] = 16'b11001_000000_00000;
        tomato_boiled[3][8] = 16'b11001_000000_00000;
        tomato_boiled[3][9] = 16'b10001_000000_00000;
        tomato_boiled[3][10] = 16'b10001_000000_00000;
        tomato_boiled[3][11] = 16'b10001_000000_00000;
        tomato_boiled[3][12] = 16'b00000_000000_00000;
        tomato_boiled[3][13] = 16'b00000_000000_00000;
        tomato_boiled[3][14] = 16'b00000_000110_11111;
        tomato_boiled[4][0] = 16'b00000_000110_11111;
        tomato_boiled[4][1] = 16'b00000_000000_00000;
        tomato_boiled[4][2] = 16'b10001_000000_00000;
        tomato_boiled[4][3] = 16'b11001_000000_00000;
        tomato_boiled[4][4] = 16'b11001_000000_00000;
        tomato_boiled[4][5] = 16'b11001_000000_00000;
        tomato_boiled[4][6] = 16'b11001_000000_00000;
        tomato_boiled[4][7] = 16'b11001_000000_00000;
        tomato_boiled[4][8] = 16'b11001_000000_00000;
        tomato_boiled[4][9] = 16'b11001_000000_00000;
        tomato_boiled[4][10] = 16'b11001_000000_00000;
        tomato_boiled[4][11] = 16'b11001_000000_00000;
        tomato_boiled[4][12] = 16'b10001_000000_00000;
        tomato_boiled[4][13] = 16'b00000_000000_00000;
        tomato_boiled[4][14] = 16'b00000_000110_11111;
        tomato_boiled[5][0] = 16'b00000_000110_11111;
        tomato_boiled[5][1] = 16'b00000_000000_00000;
        tomato_boiled[5][2] = 16'b11001_000000_00000;
        tomato_boiled[5][3] = 16'b11001_000000_00000;
        tomato_boiled[5][4] = 16'b11001_000000_00000;
        tomato_boiled[5][5] = 16'b11001_000000_00000;
        tomato_boiled[5][6] = 16'b11001_000000_00000;
        tomato_boiled[5][7] = 16'b11001_000000_00000;
        tomato_boiled[5][8] = 16'b11001_000000_00000;
        tomato_boiled[5][9] = 16'b11001_000000_00000;
        tomato_boiled[5][10] = 16'b11001_000000_00000;
        tomato_boiled[5][11] = 16'b11001_000000_00000;
        tomato_boiled[5][12] = 16'b11001_000000_00000;
        tomato_boiled[5][13] = 16'b00000_000000_00000;
        tomato_boiled[5][14] = 16'b00000_000110_11111;
        tomato_boiled[6][0] = 16'b00000_000110_11111;
        tomato_boiled[6][1] = 16'b00000_000000_00000;
        tomato_boiled[6][2] = 16'b11001_000000_00000;
        tomato_boiled[6][3] = 16'b11001_000000_00000;
        tomato_boiled[6][4] = 16'b11001_000000_00000;
        tomato_boiled[6][5] = 16'b11001_000000_00000;
        tomato_boiled[6][6] = 16'b11001_000000_00000;
        tomato_boiled[6][7] = 16'b11001_000000_00000;
        tomato_boiled[6][8] = 16'b11001_000000_00000;
        tomato_boiled[6][9] = 16'b11001_000000_00000;
        tomato_boiled[6][10] = 16'b11001_000000_00000;
        tomato_boiled[6][11] = 16'b11001_000000_00000;
        tomato_boiled[6][12] = 16'b11001_000000_00000;
        tomato_boiled[6][13] = 16'b00000_000000_00000;
        tomato_boiled[6][14] = 16'b00000_000110_11111;
        tomato_boiled[7][0] = 16'b00000_000110_11111;
        tomato_boiled[7][1] = 16'b00000_000000_00000;
        tomato_boiled[7][2] = 16'b11001_000000_00000;
        tomato_boiled[7][3] = 16'b11001_000000_00000;
        tomato_boiled[7][4] = 16'b11001_000000_00000;
        tomato_boiled[7][5] = 16'b11001_000000_00000;
        tomato_boiled[7][6] = 16'b11001_000000_00000;
        tomato_boiled[7][7] = 16'b11001_000000_00000;
        tomato_boiled[7][8] = 16'b11001_000000_00000;
        tomato_boiled[7][9] = 16'b11001_000000_00000;
        tomato_boiled[7][10] = 16'b11001_000000_00000;
        tomato_boiled[7][11] = 16'b11001_000000_00000;
        tomato_boiled[7][12] = 16'b11001_000000_00000;
        tomato_boiled[7][13] = 16'b00000_000000_00000;
        tomato_boiled[7][14] = 16'b00000_000110_11111;
        tomato_boiled[8][0] = 16'b00000_000110_11111;
        tomato_boiled[8][1] = 16'b00000_000000_00000;
        tomato_boiled[8][2] = 16'b11001_000000_00000;
        tomato_boiled[8][3] = 16'b00000_011100_00000;
        tomato_boiled[8][4] = 16'b11001_000000_00000;
        tomato_boiled[8][5] = 16'b11001_000000_00000;
        tomato_boiled[8][6] = 16'b11001_000000_00000;
        tomato_boiled[8][7] = 16'b11001_000000_00000;
        tomato_boiled[8][8] = 16'b11001_000000_00000;
        tomato_boiled[8][9] = 16'b11001_000000_00000;
        tomato_boiled[8][10] = 16'b11001_000000_00000;
        tomato_boiled[8][11] = 16'b00000_011100_00000;
        tomato_boiled[8][12] = 16'b11001_000000_00000;
        tomato_boiled[8][13] = 16'b00000_000000_00000;
        tomato_boiled[8][14] = 16'b00000_000110_11111;
        tomato_boiled[9][0] = 16'b00000_000110_11111;
        tomato_boiled[9][1] = 16'b00000_000000_00000;
        tomato_boiled[9][2] = 16'b11001_000000_00000;
        tomato_boiled[9][3] = 16'b00000_011100_00000;
        tomato_boiled[9][4] = 16'b00000_011100_00000;
        tomato_boiled[9][5] = 16'b00000_011100_00000;
        tomato_boiled[9][6] = 16'b11001_000000_00000;
        tomato_boiled[9][7] = 16'b11001_000000_00000;
        tomato_boiled[9][8] = 16'b11001_000000_00000;
        tomato_boiled[9][9] = 16'b00000_011100_00000;
        tomato_boiled[9][10] = 16'b00000_011100_00000;
        tomato_boiled[9][11] = 16'b00000_011100_00000;
        tomato_boiled[9][12] = 16'b11001_000000_00000;
        tomato_boiled[9][13] = 16'b00000_000000_00000;
        tomato_boiled[9][14] = 16'b00000_000110_11111;
        tomato_boiled[10][0] = 16'b00000_000110_11111;
        tomato_boiled[10][1] = 16'b00000_000000_00000;
        tomato_boiled[10][2] = 16'b00000_000000_00000;
        tomato_boiled[10][3] = 16'b11001_000000_00000;
        tomato_boiled[10][4] = 16'b00000_011100_00000;
        tomato_boiled[10][5] = 16'b00000_011100_00000;
        tomato_boiled[10][6] = 16'b00000_011100_00000;
        tomato_boiled[10][7] = 16'b11001_000000_00000;
        tomato_boiled[10][8] = 16'b00000_011100_00000;
        tomato_boiled[10][9] = 16'b00000_011100_00000;
        tomato_boiled[10][10] = 16'b00000_011100_00000;
        tomato_boiled[10][11] = 16'b11001_000000_00000;
        tomato_boiled[10][12] = 16'b00000_000000_00000;
        tomato_boiled[10][13] = 16'b00000_000000_00000;
        tomato_boiled[10][14] = 16'b00000_000110_11111;
        tomato_boiled[11][0] = 16'b00000_000110_11111;
        tomato_boiled[11][1] = 16'b00000_000000_00000;
        tomato_boiled[11][2] = 16'b00000_000000_00000;
        tomato_boiled[11][3] = 16'b00000_000000_00000;
        tomato_boiled[11][4] = 16'b11001_000000_00000;
        tomato_boiled[11][5] = 16'b11001_000000_00000;
        tomato_boiled[11][6] = 16'b00000_011100_00000;
        tomato_boiled[11][7] = 16'b00000_011100_00000;
        tomato_boiled[11][8] = 16'b00000_011100_00000;
        tomato_boiled[11][9] = 16'b11001_000000_00000;
        tomato_boiled[11][10] = 16'b11001_000000_00000;
        tomato_boiled[11][11] = 16'b00000_000000_00000;
        tomato_boiled[11][12] = 16'b00000_000000_00000;
        tomato_boiled[11][13] = 16'b00000_000000_00000;
        tomato_boiled[11][14] = 16'b00000_000110_11111;
        tomato_boiled[12][0] = 16'b00000_000110_11111;
        tomato_boiled[12][1] = 16'b00000_000000_00000;
        tomato_boiled[12][2] = 16'b00000_000000_00000;
        tomato_boiled[12][3] = 16'b00000_011100_00000;
        tomato_boiled[12][4] = 16'b00000_011100_00000;
        tomato_boiled[12][5] = 16'b00000_011100_00000;
        tomato_boiled[12][6] = 16'b00000_011100_00000;
        tomato_boiled[12][7] = 16'b11001_000000_00000;
        tomato_boiled[12][8] = 16'b00000_011100_00000;
        tomato_boiled[12][9] = 16'b00000_011100_00000;
        tomato_boiled[12][10] = 16'b00000_011100_00000;
        tomato_boiled[12][11] = 16'b00000_011100_00000;
        tomato_boiled[12][12] = 16'b00000_000000_00000;
        tomato_boiled[12][13] = 16'b00000_000000_00000;
        tomato_boiled[12][14] = 16'b00000_000110_11111;
        tomato_boiled[13][0] = 16'b00000_000110_11111;
        tomato_boiled[13][1] = 16'b00000_000000_00000;
        tomato_boiled[13][2] = 16'b00000_000000_00000;
        tomato_boiled[13][3] = 16'b00000_000000_00000;
        tomato_boiled[13][4] = 16'b00000_011100_00000;
        tomato_boiled[13][5] = 16'b00000_011100_00000;
        tomato_boiled[13][6] = 16'b00000_000000_00000;
        tomato_boiled[13][7] = 16'b00000_000000_00000;
        tomato_boiled[13][8] = 16'b00000_000000_00000;
        tomato_boiled[13][9] = 16'b00000_011100_00000;
        tomato_boiled[13][10] = 16'b00000_011100_00000;
        tomato_boiled[13][11] = 16'b00000_000000_00000;
        tomato_boiled[13][12] = 16'b00000_000000_00000;
        tomato_boiled[13][13] = 16'b00000_000000_00000;
        tomato_boiled[13][14] = 16'b00000_000110_11111;
        tomato_boiled[14][0] = 16'b00000_000110_11111;
        tomato_boiled[14][1] = 16'b00000_000110_11111;
        tomato_boiled[14][2] = 16'b00000_000110_11111;
        tomato_boiled[14][3] = 16'b00000_000110_11111;
        tomato_boiled[14][4] = 16'b00000_000110_11111;
        tomato_boiled[14][5] = 16'b00000_000110_11111;
        tomato_boiled[14][6] = 16'b00000_000110_11111;
        tomato_boiled[14][7] = 16'b00000_000110_11111;
        tomato_boiled[14][8] = 16'b00000_000110_11111;
        tomato_boiled[14][9] = 16'b00000_000110_11111;
        tomato_boiled[14][10] = 16'b00000_000110_11111;
        tomato_boiled[14][11] = 16'b00000_000110_11111;
        tomato_boiled[14][12] = 16'b00000_000110_11111;
        tomato_boiled[14][13] = 16'b00000_000110_11111;
        tomato_boiled[14][14] = 16'b00000_000110_11111;


        tomato_chopped[0][0] = 16'b00000_111111_00001;
        tomato_chopped[0][1] = 16'b00000_111111_00001;
        tomato_chopped[0][2] = 16'b00000_111111_00001;
        tomato_chopped[0][3] = 16'b00000_111111_00001;
        tomato_chopped[0][4] = 16'b00000_111111_00001;
        tomato_chopped[0][5] = 16'b00000_111111_00001;
        tomato_chopped[0][6] = 16'b00000_111111_00001;
        tomato_chopped[0][7] = 16'b00000_111111_00001;
        tomato_chopped[0][8] = 16'b00000_111111_00001;
        tomato_chopped[0][9] = 16'b00000_111111_00001;
        tomato_chopped[0][10] = 16'b00000_111111_00001;
        tomato_chopped[0][11] = 16'b00000_111111_00001;
        tomato_chopped[0][12] = 16'b00000_111111_00001;
        tomato_chopped[0][13] = 16'b00000_111111_00001;
        tomato_chopped[0][14] = 16'b00000_111111_00001;
        tomato_chopped[1][0] = 16'b00000_111111_00001;
        tomato_chopped[1][1] = 16'b00000_000000_00000;
        tomato_chopped[1][2] = 16'b00000_000000_00000;
        tomato_chopped[1][3] = 16'b00000_000000_00000;
        tomato_chopped[1][4] = 16'b00000_000000_00000;
        tomato_chopped[1][5] = 16'b00000_000000_00000;
        tomato_chopped[1][6] = 16'b00000_000000_00000;
        tomato_chopped[1][7] = 16'b00000_000000_00000;
        tomato_chopped[1][8] = 16'b00000_000000_00000;
        tomato_chopped[1][9] = 16'b00000_000000_00000;
        tomato_chopped[1][10] = 16'b00000_000000_00000;
        tomato_chopped[1][11] = 16'b00000_000000_00000;
        tomato_chopped[1][12] = 16'b00000_000000_00000;
        tomato_chopped[1][13] = 16'b00000_000000_00000;
        tomato_chopped[1][14] = 16'b00000_111111_00001;
        tomato_chopped[2][0] = 16'b00000_111111_00001;
        tomato_chopped[2][1] = 16'b00000_000000_00000;
        tomato_chopped[2][2] = 16'b00000_000000_00000;
        tomato_chopped[2][3] = 16'b00000_000000_00000;
        tomato_chopped[2][4] = 16'b00000_000000_00000;
        tomato_chopped[2][5] = 16'b10001_000000_00000;
        tomato_chopped[2][6] = 16'b10001_000000_00000;
        tomato_chopped[2][7] = 16'b10001_000000_00000;
        tomato_chopped[2][8] = 16'b10001_000000_00000;
        tomato_chopped[2][9] = 16'b10001_000000_00000;
        tomato_chopped[2][10] = 16'b00000_000000_00000;
        tomato_chopped[2][11] = 16'b00000_000000_00000;
        tomato_chopped[2][12] = 16'b00000_000000_00000;
        tomato_chopped[2][13] = 16'b00000_000000_00000;
        tomato_chopped[2][14] = 16'b00000_111111_00001;
        tomato_chopped[3][0] = 16'b00000_111111_00001;
        tomato_chopped[3][1] = 16'b00000_000000_00000;
        tomato_chopped[3][2] = 16'b00000_000000_00000;
        tomato_chopped[3][3] = 16'b10001_000000_00000;
        tomato_chopped[3][4] = 16'b10001_000000_00000;
        tomato_chopped[3][5] = 16'b10001_000000_00000;
        tomato_chopped[3][6] = 16'b11001_000000_00000;
        tomato_chopped[3][7] = 16'b11001_000000_00000;
        tomato_chopped[3][8] = 16'b11001_000000_00000;
        tomato_chopped[3][9] = 16'b10001_000000_00000;
        tomato_chopped[3][10] = 16'b10001_000000_00000;
        tomato_chopped[3][11] = 16'b10001_000000_00000;
        tomato_chopped[3][12] = 16'b00000_000000_00000;
        tomato_chopped[3][13] = 16'b00000_000000_00000;
        tomato_chopped[3][14] = 16'b00000_111111_00001;
        tomato_chopped[4][0] = 16'b00000_111111_00001;
        tomato_chopped[4][1] = 16'b00000_000000_00000;
        tomato_chopped[4][2] = 16'b10001_000000_00000;
        tomato_chopped[4][3] = 16'b11001_000000_00000;
        tomato_chopped[4][4] = 16'b11001_000000_00000;
        tomato_chopped[4][5] = 16'b11001_000000_00000;
        tomato_chopped[4][6] = 16'b11001_000000_00000;
        tomato_chopped[4][7] = 16'b11001_000000_00000;
        tomato_chopped[4][8] = 16'b11001_000000_00000;
        tomato_chopped[4][9] = 16'b11001_000000_00000;
        tomato_chopped[4][10] = 16'b11001_000000_00000;
        tomato_chopped[4][11] = 16'b11001_000000_00000;
        tomato_chopped[4][12] = 16'b10001_000000_00000;
        tomato_chopped[4][13] = 16'b00000_000000_00000;
        tomato_chopped[4][14] = 16'b00000_111111_00001;
        tomato_chopped[5][0] = 16'b00000_111111_00001;
        tomato_chopped[5][1] = 16'b00000_000000_00000;
        tomato_chopped[5][2] = 16'b11001_000000_00000;
        tomato_chopped[5][3] = 16'b11001_000000_00000;
        tomato_chopped[5][4] = 16'b11001_000000_00000;
        tomato_chopped[5][5] = 16'b11001_000000_00000;
        tomato_chopped[5][6] = 16'b11001_000000_00000;
        tomato_chopped[5][7] = 16'b11001_000000_00000;
        tomato_chopped[5][8] = 16'b11001_000000_00000;
        tomato_chopped[5][9] = 16'b11001_000000_00000;
        tomato_chopped[5][10] = 16'b11001_000000_00000;
        tomato_chopped[5][11] = 16'b11001_000000_00000;
        tomato_chopped[5][12] = 16'b11001_000000_00000;
        tomato_chopped[5][13] = 16'b00000_000000_00000;
        tomato_chopped[5][14] = 16'b00000_111111_00001;
        tomato_chopped[6][0] = 16'b00000_111111_00001;
        tomato_chopped[6][1] = 16'b00000_000000_00000;
        tomato_chopped[6][2] = 16'b11001_000000_00000;
        tomato_chopped[6][3] = 16'b11001_000000_00000;
        tomato_chopped[6][4] = 16'b11001_000000_00000;
        tomato_chopped[6][5] = 16'b11001_000000_00000;
        tomato_chopped[6][6] = 16'b11001_000000_00000;
        tomato_chopped[6][7] = 16'b11001_000000_00000;
        tomato_chopped[6][8] = 16'b11001_000000_00000;
        tomato_chopped[6][9] = 16'b11001_000000_00000;
        tomato_chopped[6][10] = 16'b11001_000000_00000;
        tomato_chopped[6][11] = 16'b11001_000000_00000;
        tomato_chopped[6][12] = 16'b11001_000000_00000;
        tomato_chopped[6][13] = 16'b00000_000000_00000;
        tomato_chopped[6][14] = 16'b00000_111111_00001;
        tomato_chopped[7][0] = 16'b00000_111111_00001;
        tomato_chopped[7][1] = 16'b00000_000000_00000;
        tomato_chopped[7][2] = 16'b11001_000000_00000;
        tomato_chopped[7][3] = 16'b11001_000000_00000;
        tomato_chopped[7][4] = 16'b11001_000000_00000;
        tomato_chopped[7][5] = 16'b11001_000000_00000;
        tomato_chopped[7][6] = 16'b11001_000000_00000;
        tomato_chopped[7][7] = 16'b11001_000000_00000;
        tomato_chopped[7][8] = 16'b11001_000000_00000;
        tomato_chopped[7][9] = 16'b11001_000000_00000;
        tomato_chopped[7][10] = 16'b11001_000000_00000;
        tomato_chopped[7][11] = 16'b11001_000000_00000;
        tomato_chopped[7][12] = 16'b11001_000000_00000;
        tomato_chopped[7][13] = 16'b00000_000000_00000;
        tomato_chopped[7][14] = 16'b00000_111111_00001;
        tomato_chopped[8][0] = 16'b00000_111111_00001;
        tomato_chopped[8][1] = 16'b00000_000000_00000;
        tomato_chopped[8][2] = 16'b11001_000000_00000;
        tomato_chopped[8][3] = 16'b00000_011100_00000;
        tomato_chopped[8][4] = 16'b11001_000000_00000;
        tomato_chopped[8][5] = 16'b11001_000000_00000;
        tomato_chopped[8][6] = 16'b11001_000000_00000;
        tomato_chopped[8][7] = 16'b11001_000000_00000;
        tomato_chopped[8][8] = 16'b11001_000000_00000;
        tomato_chopped[8][9] = 16'b11001_000000_00000;
        tomato_chopped[8][10] = 16'b11001_000000_00000;
        tomato_chopped[8][11] = 16'b00000_011100_00000;
        tomato_chopped[8][12] = 16'b11001_000000_00000;
        tomato_chopped[8][13] = 16'b00000_000000_00000;
        tomato_chopped[8][14] = 16'b00000_111111_00001;
        tomato_chopped[9][0] = 16'b00000_111111_00001;
        tomato_chopped[9][1] = 16'b00000_000000_00000;
        tomato_chopped[9][2] = 16'b11001_000000_00000;
        tomato_chopped[9][3] = 16'b00000_011100_00000;
        tomato_chopped[9][4] = 16'b00000_011100_00000;
        tomato_chopped[9][5] = 16'b00000_011100_00000;
        tomato_chopped[9][6] = 16'b11001_000000_00000;
        tomato_chopped[9][7] = 16'b11001_000000_00000;
        tomato_chopped[9][8] = 16'b11001_000000_00000;
        tomato_chopped[9][9] = 16'b00000_011100_00000;
        tomato_chopped[9][10] = 16'b00000_011100_00000;
        tomato_chopped[9][11] = 16'b00000_011100_00000;
        tomato_chopped[9][12] = 16'b11001_000000_00000;
        tomato_chopped[9][13] = 16'b00000_000000_00000;
        tomato_chopped[9][14] = 16'b00000_111111_00001;
        tomato_chopped[10][0] = 16'b00000_111111_00001;
        tomato_chopped[10][1] = 16'b00000_000000_00000;
        tomato_chopped[10][2] = 16'b00000_000000_00000;
        tomato_chopped[10][3] = 16'b11001_000000_00000;
        tomato_chopped[10][4] = 16'b00000_011100_00000;
        tomato_chopped[10][5] = 16'b00000_011100_00000;
        tomato_chopped[10][6] = 16'b00000_011100_00000;
        tomato_chopped[10][7] = 16'b11001_000000_00000;
        tomato_chopped[10][8] = 16'b00000_011100_00000;
        tomato_chopped[10][9] = 16'b00000_011100_00000;
        tomato_chopped[10][10] = 16'b00000_011100_00000;
        tomato_chopped[10][11] = 16'b11001_000000_00000;
        tomato_chopped[10][12] = 16'b00000_000000_00000;
        tomato_chopped[10][13] = 16'b00000_000000_00000;
        tomato_chopped[10][14] = 16'b00000_111111_00001;
        tomato_chopped[11][0] = 16'b00000_111111_00001;
        tomato_chopped[11][1] = 16'b00000_000000_00000;
        tomato_chopped[11][2] = 16'b00000_000000_00000;
        tomato_chopped[11][3] = 16'b00000_000000_00000;
        tomato_chopped[11][4] = 16'b11001_000000_00000;
        tomato_chopped[11][5] = 16'b11001_000000_00000;
        tomato_chopped[11][6] = 16'b00000_011100_00000;
        tomato_chopped[11][7] = 16'b00000_011100_00000;
        tomato_chopped[11][8] = 16'b00000_011100_00000;
        tomato_chopped[11][9] = 16'b11001_000000_00000;
        tomato_chopped[11][10] = 16'b11001_000000_00000;
        tomato_chopped[11][11] = 16'b00000_000000_00000;
        tomato_chopped[11][12] = 16'b00000_000000_00000;
        tomato_chopped[11][13] = 16'b00000_000000_00000;
        tomato_chopped[11][14] = 16'b00000_111111_00001;
        tomato_chopped[12][0] = 16'b00000_111111_00001;
        tomato_chopped[12][1] = 16'b00000_000000_00000;
        tomato_chopped[12][2] = 16'b00000_000000_00000;
        tomato_chopped[12][3] = 16'b00000_011100_00000;
        tomato_chopped[12][4] = 16'b00000_011100_00000;
        tomato_chopped[12][5] = 16'b00000_011100_00000;
        tomato_chopped[12][6] = 16'b00000_011100_00000;
        tomato_chopped[12][7] = 16'b11001_000000_00000;
        tomato_chopped[12][8] = 16'b00000_011100_00000;
        tomato_chopped[12][9] = 16'b00000_011100_00000;
        tomato_chopped[12][10] = 16'b00000_011100_00000;
        tomato_chopped[12][11] = 16'b00000_011100_00000;
        tomato_chopped[12][12] = 16'b00000_000000_00000;
        tomato_chopped[12][13] = 16'b00000_000000_00000;
        tomato_chopped[12][14] = 16'b00000_111111_00001;
        tomato_chopped[13][0] = 16'b00000_111111_00001;
        tomato_chopped[13][1] = 16'b00000_000000_00000;
        tomato_chopped[13][2] = 16'b00000_000000_00000;
        tomato_chopped[13][3] = 16'b00000_000000_00000;
        tomato_chopped[13][4] = 16'b00000_011100_00000;
        tomato_chopped[13][5] = 16'b00000_011100_00000;
        tomato_chopped[13][6] = 16'b00000_000000_00000;
        tomato_chopped[13][7] = 16'b00000_000000_00000;
        tomato_chopped[13][8] = 16'b00000_000000_00000;
        tomato_chopped[13][9] = 16'b00000_011100_00000;
        tomato_chopped[13][10] = 16'b00000_011100_00000;
        tomato_chopped[13][11] = 16'b00000_000000_00000;
        tomato_chopped[13][12] = 16'b00000_000000_00000;
        tomato_chopped[13][13] = 16'b00000_000000_00000;
        tomato_chopped[13][14] = 16'b00000_111111_00001;
        tomato_chopped[14][0] = 16'b00000_111111_00001;
        tomato_chopped[14][1] = 16'b00000_111111_00001;
        tomato_chopped[14][2] = 16'b00000_111111_00001;
        tomato_chopped[14][3] = 16'b00000_111111_00001;
        tomato_chopped[14][4] = 16'b00000_111111_00001;
        tomato_chopped[14][5] = 16'b00000_111111_00001;
        tomato_chopped[14][6] = 16'b00000_111111_00001;
        tomato_chopped[14][7] = 16'b00000_111111_00001;
        tomato_chopped[14][8] = 16'b00000_111111_00001;
        tomato_chopped[14][9] = 16'b00000_111111_00001;
        tomato_chopped[14][10] = 16'b00000_111111_00001;
        tomato_chopped[14][11] = 16'b00000_111111_00001;
        tomato_chopped[14][12] = 16'b00000_111111_00001;
        tomato_chopped[14][13] = 16'b00000_111111_00001;
        tomato_chopped[14][14] = 16'b00000_111111_00001;


        tomato_raw[0][0] = 16'b11001_000000_00000;
        tomato_raw[0][1] = 16'b11001_000000_00000;
        tomato_raw[0][2] = 16'b11001_000000_00000;
        tomato_raw[0][3] = 16'b11001_000000_00000;
        tomato_raw[0][4] = 16'b11001_000000_00000;
        tomato_raw[0][5] = 16'b11001_000000_00000;
        tomato_raw[0][6] = 16'b11001_000000_00000;
        tomato_raw[0][7] = 16'b11001_000000_00000;
        tomato_raw[0][8] = 16'b11001_000000_00000;
        tomato_raw[0][9] = 16'b11001_000000_00000;
        tomato_raw[0][10] = 16'b11001_000000_00000;
        tomato_raw[0][11] = 16'b11001_000000_00000;
        tomato_raw[0][12] = 16'b11001_000000_00000;
        tomato_raw[0][13] = 16'b11001_000000_00000;
        tomato_raw[0][14] = 16'b11001_000000_00000;
        tomato_raw[1][0] = 16'b11001_000000_00000;
        tomato_raw[1][1] = 16'b00000_000000_00000;
        tomato_raw[1][2] = 16'b00000_000000_00000;
        tomato_raw[1][3] = 16'b00000_000000_00000;
        tomato_raw[1][4] = 16'b00000_000000_00000;
        tomato_raw[1][5] = 16'b00000_000000_00000;
        tomato_raw[1][6] = 16'b00000_000000_00000;
        tomato_raw[1][7] = 16'b00000_000000_00000;
        tomato_raw[1][8] = 16'b00000_000000_00000;
        tomato_raw[1][9] = 16'b00000_000000_00000;
        tomato_raw[1][10] = 16'b00000_000000_00000;
        tomato_raw[1][11] = 16'b00000_000000_00000;
        tomato_raw[1][12] = 16'b00000_000000_00000;
        tomato_raw[1][13] = 16'b00000_000000_00000;
        tomato_raw[1][14] = 16'b11001_000000_00000;
        tomato_raw[2][0] = 16'b11001_000000_00000;
        tomato_raw[2][1] = 16'b00000_000000_00000;
        tomato_raw[2][2] = 16'b00000_000000_00000;
        tomato_raw[2][3] = 16'b00000_000000_00000;
        tomato_raw[2][4] = 16'b00000_000000_00000;
        tomato_raw[2][5] = 16'b10001_000000_00000;
        tomato_raw[2][6] = 16'b10001_000000_00000;
        tomato_raw[2][7] = 16'b10001_000000_00000;
        tomato_raw[2][8] = 16'b10001_000000_00000;
        tomato_raw[2][9] = 16'b10001_000000_00000;
        tomato_raw[2][10] = 16'b00000_000000_00000;
        tomato_raw[2][11] = 16'b00000_000000_00000;
        tomato_raw[2][12] = 16'b00000_000000_00000;
        tomato_raw[2][13] = 16'b00000_000000_00000;
        tomato_raw[2][14] = 16'b11001_000000_00000;
        tomato_raw[3][0] = 16'b11001_000000_00000;
        tomato_raw[3][1] = 16'b00000_000000_00000;
        tomato_raw[3][2] = 16'b00000_000000_00000;
        tomato_raw[3][3] = 16'b10001_000000_00000;
        tomato_raw[3][4] = 16'b10001_000000_00000;
        tomato_raw[3][5] = 16'b10001_000000_00000;
        tomato_raw[3][6] = 16'b11001_000000_00000;
        tomato_raw[3][7] = 16'b11001_000000_00000;
        tomato_raw[3][8] = 16'b11001_000000_00000;
        tomato_raw[3][9] = 16'b10001_000000_00000;
        tomato_raw[3][10] = 16'b10001_000000_00000;
        tomato_raw[3][11] = 16'b10001_000000_00000;
        tomato_raw[3][12] = 16'b00000_000000_00000;
        tomato_raw[3][13] = 16'b00000_000000_00000;
        tomato_raw[3][14] = 16'b11001_000000_00000;
        tomato_raw[4][0] = 16'b11001_000000_00000;
        tomato_raw[4][1] = 16'b00000_000000_00000;
        tomato_raw[4][2] = 16'b10001_000000_00000;
        tomato_raw[4][3] = 16'b11001_000000_00000;
        tomato_raw[4][4] = 16'b11001_000000_00000;
        tomato_raw[4][5] = 16'b11001_000000_00000;
        tomato_raw[4][6] = 16'b11001_000000_00000;
        tomato_raw[4][7] = 16'b11001_000000_00000;
        tomato_raw[4][8] = 16'b11001_000000_00000;
        tomato_raw[4][9] = 16'b11001_000000_00000;
        tomato_raw[4][10] = 16'b11001_000000_00000;
        tomato_raw[4][11] = 16'b11001_000000_00000;
        tomato_raw[4][12] = 16'b10001_000000_00000;
        tomato_raw[4][13] = 16'b00000_000000_00000;
        tomato_raw[4][14] = 16'b11001_000000_00000;
        tomato_raw[5][0] = 16'b11001_000000_00000;
        tomato_raw[5][1] = 16'b00000_000000_00000;
        tomato_raw[5][2] = 16'b11001_000000_00000;
        tomato_raw[5][3] = 16'b11001_000000_00000;
        tomato_raw[5][4] = 16'b11001_000000_00000;
        tomato_raw[5][5] = 16'b11001_000000_00000;
        tomato_raw[5][6] = 16'b11001_000000_00000;
        tomato_raw[5][7] = 16'b11001_000000_00000;
        tomato_raw[5][8] = 16'b11001_000000_00000;
        tomato_raw[5][9] = 16'b11001_000000_00000;
        tomato_raw[5][10] = 16'b11001_000000_00000;
        tomato_raw[5][11] = 16'b11001_000000_00000;
        tomato_raw[5][12] = 16'b11001_000000_00000;
        tomato_raw[5][13] = 16'b00000_000000_00000;
        tomato_raw[5][14] = 16'b11001_000000_00000;
        tomato_raw[6][0] = 16'b11001_000000_00000;
        tomato_raw[6][1] = 16'b00000_000000_00000;
        tomato_raw[6][2] = 16'b11001_000000_00000;
        tomato_raw[6][3] = 16'b11001_000000_00000;
        tomato_raw[6][4] = 16'b11001_000000_00000;
        tomato_raw[6][5] = 16'b11001_000000_00000;
        tomato_raw[6][6] = 16'b11001_000000_00000;
        tomato_raw[6][7] = 16'b11001_000000_00000;
        tomato_raw[6][8] = 16'b11001_000000_00000;
        tomato_raw[6][9] = 16'b11001_000000_00000;
        tomato_raw[6][10] = 16'b11001_000000_00000;
        tomato_raw[6][11] = 16'b11001_000000_00000;
        tomato_raw[6][12] = 16'b11001_000000_00000;
        tomato_raw[6][13] = 16'b00000_000000_00000;
        tomato_raw[6][14] = 16'b11001_000000_00000;
        tomato_raw[7][0] = 16'b11001_000000_00000;
        tomato_raw[7][1] = 16'b00000_000000_00000;
        tomato_raw[7][2] = 16'b11001_000000_00000;
        tomato_raw[7][3] = 16'b11001_000000_00000;
        tomato_raw[7][4] = 16'b11001_000000_00000;
        tomato_raw[7][5] = 16'b11001_000000_00000;
        tomato_raw[7][6] = 16'b11001_000000_00000;
        tomato_raw[7][7] = 16'b11001_000000_00000;
        tomato_raw[7][8] = 16'b11001_000000_00000;
        tomato_raw[7][9] = 16'b11001_000000_00000;
        tomato_raw[7][10] = 16'b11001_000000_00000;
        tomato_raw[7][11] = 16'b11001_000000_00000;
        tomato_raw[7][12] = 16'b11001_000000_00000;
        tomato_raw[7][13] = 16'b00000_000000_00000;
        tomato_raw[7][14] = 16'b11001_000000_00000;
        tomato_raw[8][0] = 16'b11001_000000_00000;
        tomato_raw[8][1] = 16'b00000_000000_00000;
        tomato_raw[8][2] = 16'b11001_000000_00000;
        tomato_raw[8][3] = 16'b00000_011100_00000;
        tomato_raw[8][4] = 16'b11001_000000_00000;
        tomato_raw[8][5] = 16'b11001_000000_00000;
        tomato_raw[8][6] = 16'b11001_000000_00000;
        tomato_raw[8][7] = 16'b11001_000000_00000;
        tomato_raw[8][8] = 16'b11001_000000_00000;
        tomato_raw[8][9] = 16'b11001_000000_00000;
        tomato_raw[8][10] = 16'b11001_000000_00000;
        tomato_raw[8][11] = 16'b00000_011100_00000;
        tomato_raw[8][12] = 16'b11001_000000_00000;
        tomato_raw[8][13] = 16'b00000_000000_00000;
        tomato_raw[8][14] = 16'b11001_000000_00000;
        tomato_raw[9][0] = 16'b11001_000000_00000;
        tomato_raw[9][1] = 16'b00000_000000_00000;
        tomato_raw[9][2] = 16'b11001_000000_00000;
        tomato_raw[9][3] = 16'b00000_011100_00000;
        tomato_raw[9][4] = 16'b00000_011100_00000;
        tomato_raw[9][5] = 16'b00000_011100_00000;
        tomato_raw[9][6] = 16'b11001_000000_00000;
        tomato_raw[9][7] = 16'b11001_000000_00000;
        tomato_raw[9][8] = 16'b11001_000000_00000;
        tomato_raw[9][9] = 16'b00000_011100_00000;
        tomato_raw[9][10] = 16'b00000_011100_00000;
        tomato_raw[9][11] = 16'b00000_011100_00000;
        tomato_raw[9][12] = 16'b11001_000000_00000;
        tomato_raw[9][13] = 16'b00000_000000_00000;
        tomato_raw[9][14] = 16'b11001_000000_00000;
        tomato_raw[10][0] = 16'b11001_000000_00000;
        tomato_raw[10][1] = 16'b00000_000000_00000;
        tomato_raw[10][2] = 16'b00000_000000_00000;
        tomato_raw[10][3] = 16'b11001_000000_00000;
        tomato_raw[10][4] = 16'b00000_011100_00000;
        tomato_raw[10][5] = 16'b00000_011100_00000;
        tomato_raw[10][6] = 16'b00000_011100_00000;
        tomato_raw[10][7] = 16'b11001_000000_00000;
        tomato_raw[10][8] = 16'b00000_011100_00000;
        tomato_raw[10][9] = 16'b00000_011100_00000;
        tomato_raw[10][10] = 16'b00000_011100_00000;
        tomato_raw[10][11] = 16'b11001_000000_00000;
        tomato_raw[10][12] = 16'b00000_000000_00000;
        tomato_raw[10][13] = 16'b00000_000000_00000;
        tomato_raw[10][14] = 16'b11001_000000_00000;
        tomato_raw[11][0] = 16'b11001_000000_00000;
        tomato_raw[11][1] = 16'b00000_000000_00000;
        tomato_raw[11][2] = 16'b00000_000000_00000;
        tomato_raw[11][3] = 16'b00000_000000_00000;
        tomato_raw[11][4] = 16'b11001_000000_00000;
        tomato_raw[11][5] = 16'b11001_000000_00000;
        tomato_raw[11][6] = 16'b00000_011100_00000;
        tomato_raw[11][7] = 16'b00000_011100_00000;
        tomato_raw[11][8] = 16'b00000_011100_00000;
        tomato_raw[11][9] = 16'b11001_000000_00000;
        tomato_raw[11][10] = 16'b11001_000000_00000;
        tomato_raw[11][11] = 16'b00000_000000_00000;
        tomato_raw[11][12] = 16'b00000_000000_00000;
        tomato_raw[11][13] = 16'b00000_000000_00000;
        tomato_raw[11][14] = 16'b11001_000000_00000;
        tomato_raw[12][0] = 16'b11001_000000_00000;
        tomato_raw[12][1] = 16'b00000_000000_00000;
        tomato_raw[12][2] = 16'b00000_000000_00000;
        tomato_raw[12][3] = 16'b00000_011100_00000;
        tomato_raw[12][4] = 16'b00000_011100_00000;
        tomato_raw[12][5] = 16'b00000_011100_00000;
        tomato_raw[12][6] = 16'b00000_011100_00000;
        tomato_raw[12][7] = 16'b11001_000000_00000;
        tomato_raw[12][8] = 16'b00000_011100_00000;
        tomato_raw[12][9] = 16'b00000_011100_00000;
        tomato_raw[12][10] = 16'b00000_011100_00000;
        tomato_raw[12][11] = 16'b00000_011100_00000;
        tomato_raw[12][12] = 16'b00000_000000_00000;
        tomato_raw[12][13] = 16'b00000_000000_00000;
        tomato_raw[12][14] = 16'b11001_000000_00000;
        tomato_raw[13][0] = 16'b11001_000000_00000;
        tomato_raw[13][1] = 16'b00000_000000_00000;
        tomato_raw[13][2] = 16'b00000_000000_00000;
        tomato_raw[13][3] = 16'b00000_000000_00000;
        tomato_raw[13][4] = 16'b00000_011100_00000;
        tomato_raw[13][5] = 16'b00000_011100_00000;
        tomato_raw[13][6] = 16'b00000_000000_00000;
        tomato_raw[13][7] = 16'b00000_000000_00000;
        tomato_raw[13][8] = 16'b00000_000000_00000;
        tomato_raw[13][9] = 16'b00000_011100_00000;
        tomato_raw[13][10] = 16'b00000_011100_00000;
        tomato_raw[13][11] = 16'b00000_000000_00000;
        tomato_raw[13][12] = 16'b00000_000000_00000;
        tomato_raw[13][13] = 16'b00000_000000_00000;
        tomato_raw[13][14] = 16'b11001_000000_00000;
        tomato_raw[14][0] = 16'b11001_000000_00000;
        tomato_raw[14][1] = 16'b11001_000000_00000;
        tomato_raw[14][2] = 16'b11001_000000_00000;
        tomato_raw[14][3] = 16'b11001_000000_00000;
        tomato_raw[14][4] = 16'b11001_000000_00000;
        tomato_raw[14][5] = 16'b11001_000000_00000;
        tomato_raw[14][6] = 16'b11001_000000_00000;
        tomato_raw[14][7] = 16'b11001_000000_00000;
        tomato_raw[14][8] = 16'b11001_000000_00000;
        tomato_raw[14][9] = 16'b11001_000000_00000;
        tomato_raw[14][10] = 16'b11001_000000_00000;
        tomato_raw[14][11] = 16'b11001_000000_00000;
        tomato_raw[14][12] = 16'b11001_000000_00000;
        tomato_raw[14][13] = 16'b11001_000000_00000;
        tomato_raw[14][14] = 16'b11001_000000_00000;
        
        
        tick_overlay[0][0] = 16'b00000_101101_00000;
        tick_overlay[0][1] = 16'b00000_101101_00000;
        tick_overlay[0][2] = 16'b00000_101101_00000;
        tick_overlay[0][3] = 16'b00000_101101_00000;
        tick_overlay[0][4] = 16'b00000_101101_00000;
        tick_overlay[0][5] = 16'b00000_101101_00000;
        tick_overlay[0][6] = 16'b00000_101101_00000;
        tick_overlay[0][7] = 16'b00000_101101_00000;
        tick_overlay[0][8] = 16'b00000_101101_00000;
        tick_overlay[0][9] = 16'b00000_101101_00000;
        tick_overlay[0][10] = 16'b00000_101101_00000;
        tick_overlay[0][11] = 16'b00000_101101_00000;
        tick_overlay[0][12] = 16'b00000_101101_00000;
        tick_overlay[0][13] = 16'b00000_101101_00000;
        tick_overlay[0][14] = 16'b00000_101101_00000;
        tick_overlay[0][15] = 16'b00000_101101_00000;
        tick_overlay[0][16] = 16'b00000_101101_00000;
        tick_overlay[0][17] = 16'b00000_101101_00000;
        tick_overlay[0][18] = 16'b00000_101101_00000;
        tick_overlay[0][19] = 16'b00000_101101_00000;
        tick_overlay[0][20] = 16'b00000_101101_00000;
        tick_overlay[0][21] = 16'b00000_101101_00000;
        tick_overlay[0][22] = 16'b00000_101101_00000;
        tick_overlay[0][23] = 16'b00000_101101_00000;
        tick_overlay[0][24] = 16'b00000_101101_00000;
        tick_overlay[0][25] = 16'b00000_101101_00000;
        tick_overlay[0][26] = 16'b00000_101101_00000;
        tick_overlay[0][27] = 16'b00000_101101_00000;
        tick_overlay[0][28] = 16'b00000_101101_00000;
        tick_overlay[0][29] = 16'b00000_101101_00000;
        tick_overlay[0][30] = 16'b00000_101101_00000;
        tick_overlay[0][31] = 16'b00000_101101_00000;
        tick_overlay[1][0] = 16'b00000_101101_00000;
        tick_overlay[1][1] = 16'b00000_101101_00000;
        tick_overlay[1][2] = 16'b00000_101101_00000;
        tick_overlay[1][3] = 16'b00000_101101_00000;
        tick_overlay[1][4] = 16'b00000_101101_00000;
        tick_overlay[1][5] = 16'b00000_101101_00000;
        tick_overlay[1][6] = 16'b00000_101101_00000;
        tick_overlay[1][7] = 16'b00000_101101_00000;
        tick_overlay[1][8] = 16'b00000_101101_00000;
        tick_overlay[1][9] = 16'b00000_101101_00000;
        tick_overlay[1][10] = 16'b00000_101101_00000;
        tick_overlay[1][11] = 16'b00000_101101_00000;
        tick_overlay[1][12] = 16'b00000_101101_00000;
        tick_overlay[1][13] = 16'b00000_101101_00000;
        tick_overlay[1][14] = 16'b00000_101101_00000;
        tick_overlay[1][15] = 16'b00000_101101_00000;
        tick_overlay[1][16] = 16'b00000_101101_00000;
        tick_overlay[1][17] = 16'b00000_101101_00000;
        tick_overlay[1][18] = 16'b00000_101101_00000;
        tick_overlay[1][19] = 16'b00000_101101_00000;
        tick_overlay[1][20] = 16'b00000_101101_00000;
        tick_overlay[1][21] = 16'b00000_101101_00000;
        tick_overlay[1][22] = 16'b00000_101101_00000;
        tick_overlay[1][23] = 16'b00000_101101_00000;
        tick_overlay[1][24] = 16'b00000_101101_00000;
        tick_overlay[1][25] = 16'b00000_101101_00000;
        tick_overlay[1][26] = 16'b00000_101101_00000;
        tick_overlay[1][27] = 16'b00000_101101_00000;
        tick_overlay[1][28] = 16'b00000_101101_00000;
        tick_overlay[1][29] = 16'b00000_101101_00000;
        tick_overlay[1][30] = 16'b00000_101101_00000;
        tick_overlay[1][31] = 16'b00000_101101_00000;
        tick_overlay[2][0] = 16'b00000_101101_00000;
        tick_overlay[2][1] = 16'b00000_101101_00000;
        tick_overlay[2][2] = 16'b00000_000000_00000;
        tick_overlay[2][3] = 16'b00000_000000_00000;
        tick_overlay[2][4] = 16'b00000_000000_00000;
        tick_overlay[2][5] = 16'b00000_000000_00000;
        tick_overlay[2][6] = 16'b00000_000000_00000;
        tick_overlay[2][7] = 16'b00000_000000_00000;
        tick_overlay[2][8] = 16'b00000_000000_00000;
        tick_overlay[2][9] = 16'b00000_000000_00000;
        tick_overlay[2][10] = 16'b00000_000000_00000;
        tick_overlay[2][11] = 16'b00000_000000_00000;
        tick_overlay[2][12] = 16'b00000_000000_00000;
        tick_overlay[2][13] = 16'b00000_000000_00000;
        tick_overlay[2][14] = 16'b00000_000000_00000;
        tick_overlay[2][15] = 16'b00000_000000_00000;
        tick_overlay[2][16] = 16'b00000_000000_00000;
        tick_overlay[2][17] = 16'b00000_000000_00000;
        tick_overlay[2][18] = 16'b00000_000000_00000;
        tick_overlay[2][19] = 16'b00000_000000_00000;
        tick_overlay[2][20] = 16'b00000_000000_00000;
        tick_overlay[2][21] = 16'b00000_000000_00000;
        tick_overlay[2][22] = 16'b00000_000000_00000;
        tick_overlay[2][23] = 16'b00000_000000_00000;
        tick_overlay[2][24] = 16'b00000_000000_00000;
        tick_overlay[2][25] = 16'b00000_000000_00000;
        tick_overlay[2][26] = 16'b00000_000000_00000;
        tick_overlay[2][27] = 16'b00000_000000_00000;
        tick_overlay[2][28] = 16'b00000_000000_00000;
        tick_overlay[2][29] = 16'b00000_000000_00000;
        tick_overlay[2][30] = 16'b00000_101101_00000;
        tick_overlay[2][31] = 16'b00000_101101_00000;
        tick_overlay[3][0] = 16'b00000_101101_00000;
        tick_overlay[3][1] = 16'b00000_101101_00000;
        tick_overlay[3][2] = 16'b00000_000000_00000;
        tick_overlay[3][3] = 16'b00000_000000_00000;
        tick_overlay[3][4] = 16'b00000_000000_00000;
        tick_overlay[3][5] = 16'b00000_000000_00000;
        tick_overlay[3][6] = 16'b00000_000000_00000;
        tick_overlay[3][7] = 16'b00000_000000_00000;
        tick_overlay[3][8] = 16'b00000_000000_00000;
        tick_overlay[3][9] = 16'b00000_000000_00000;
        tick_overlay[3][10] = 16'b00000_000000_00000;
        tick_overlay[3][11] = 16'b00000_000000_00000;
        tick_overlay[3][12] = 16'b00000_000000_00000;
        tick_overlay[3][13] = 16'b00000_000000_00000;
        tick_overlay[3][14] = 16'b00000_000000_00000;
        tick_overlay[3][15] = 16'b00000_000000_00000;
        tick_overlay[3][16] = 16'b00000_000000_00000;
        tick_overlay[3][17] = 16'b00000_000000_00000;
        tick_overlay[3][18] = 16'b00000_000000_00000;
        tick_overlay[3][19] = 16'b00000_000000_00000;
        tick_overlay[3][20] = 16'b00000_000000_00000;
        tick_overlay[3][21] = 16'b00000_000000_00000;
        tick_overlay[3][22] = 16'b00000_000000_00000;
        tick_overlay[3][23] = 16'b00000_000000_00000;
        tick_overlay[3][24] = 16'b00000_000000_00000;
        tick_overlay[3][25] = 16'b00000_000000_00000;
        tick_overlay[3][26] = 16'b00000_000000_00000;
        tick_overlay[3][27] = 16'b00000_000000_00000;
        tick_overlay[3][28] = 16'b00000_000000_00000;
        tick_overlay[3][29] = 16'b00000_000000_00000;
        tick_overlay[3][30] = 16'b00000_101101_00000;
        tick_overlay[3][31] = 16'b00000_101101_00000;
        tick_overlay[4][0] = 16'b00000_101101_00000;
        tick_overlay[4][1] = 16'b00000_101101_00000;
        tick_overlay[4][2] = 16'b00000_000000_00000;
        tick_overlay[4][3] = 16'b00000_000000_00000;
        tick_overlay[4][4] = 16'b00000_000000_00000;
        tick_overlay[4][5] = 16'b00000_000000_00000;
        tick_overlay[4][6] = 16'b00000_000000_00000;
        tick_overlay[4][7] = 16'b00000_000000_00000;
        tick_overlay[4][8] = 16'b00000_000000_00000;
        tick_overlay[4][9] = 16'b00000_000000_00000;
        tick_overlay[4][10] = 16'b00000_000000_00000;
        tick_overlay[4][11] = 16'b00000_000000_00000;
        tick_overlay[4][12] = 16'b00000_000000_00000;
        tick_overlay[4][13] = 16'b00000_000000_00000;
        tick_overlay[4][14] = 16'b00000_000000_00000;
        tick_overlay[4][15] = 16'b00000_000000_00000;
        tick_overlay[4][16] = 16'b00000_000000_00000;
        tick_overlay[4][17] = 16'b00000_000000_00000;
        tick_overlay[4][18] = 16'b00000_000000_00000;
        tick_overlay[4][19] = 16'b00000_000000_00000;
        tick_overlay[4][20] = 16'b00000_000000_00000;
        tick_overlay[4][21] = 16'b00000_000000_00000;
        tick_overlay[4][22] = 16'b00000_000000_00000;
        tick_overlay[4][23] = 16'b00000_000000_00000;
        tick_overlay[4][24] = 16'b00000_000000_00000;
        tick_overlay[4][25] = 16'b00000_000000_00000;
        tick_overlay[4][26] = 16'b00000_000000_00000;
        tick_overlay[4][27] = 16'b00000_000000_00000;
        tick_overlay[4][28] = 16'b00000_000000_00000;
        tick_overlay[4][29] = 16'b00000_000000_00000;
        tick_overlay[4][30] = 16'b00000_101101_00000;
        tick_overlay[4][31] = 16'b00000_101101_00000;
        tick_overlay[5][0] = 16'b00000_101101_00000;
        tick_overlay[5][1] = 16'b00000_101101_00000;
        tick_overlay[5][2] = 16'b00000_000000_00000;
        tick_overlay[5][3] = 16'b00000_000000_00000;
        tick_overlay[5][4] = 16'b00000_000000_00000;
        tick_overlay[5][5] = 16'b00000_000000_00000;
        tick_overlay[5][6] = 16'b00000_000000_00000;
        tick_overlay[5][7] = 16'b00000_000000_00000;
        tick_overlay[5][8] = 16'b00000_000000_00000;
        tick_overlay[5][9] = 16'b00000_000000_00000;
        tick_overlay[5][10] = 16'b00000_000000_00000;
        tick_overlay[5][11] = 16'b00000_000000_00000;
        tick_overlay[5][12] = 16'b00000_000000_00000;
        tick_overlay[5][13] = 16'b00000_000000_00000;
        tick_overlay[5][14] = 16'b00000_000000_00000;
        tick_overlay[5][15] = 16'b00000_000000_00000;
        tick_overlay[5][16] = 16'b00000_000000_00000;
        tick_overlay[5][17] = 16'b00000_000000_00000;
        tick_overlay[5][18] = 16'b00000_000000_00000;
        tick_overlay[5][19] = 16'b00000_000000_00000;
        tick_overlay[5][20] = 16'b00000_000000_00000;
        tick_overlay[5][21] = 16'b00000_000000_00000;
        tick_overlay[5][22] = 16'b00000_000000_00000;
        tick_overlay[5][23] = 16'b00000_000000_00000;
        tick_overlay[5][24] = 16'b00000_000000_00000;
        tick_overlay[5][25] = 16'b00000_000000_00000;
        tick_overlay[5][26] = 16'b00000_000000_00000;
        tick_overlay[5][27] = 16'b00000_000000_00000;
        tick_overlay[5][28] = 16'b00000_000000_00000;
        tick_overlay[5][29] = 16'b00000_000000_00000;
        tick_overlay[5][30] = 16'b00000_101101_00000;
        tick_overlay[5][31] = 16'b00000_101101_00000;
        tick_overlay[6][0] = 16'b00000_101101_00000;
        tick_overlay[6][1] = 16'b00000_101101_00000;
        tick_overlay[6][2] = 16'b00000_000000_00000;
        tick_overlay[6][3] = 16'b00000_000000_00000;
        tick_overlay[6][4] = 16'b00000_000000_00000;
        tick_overlay[6][5] = 16'b00000_000000_00000;
        tick_overlay[6][6] = 16'b00000_000000_00000;
        tick_overlay[6][7] = 16'b00000_000000_00000;
        tick_overlay[6][8] = 16'b00000_000000_00000;
        tick_overlay[6][9] = 16'b00000_000000_00000;
        tick_overlay[6][10] = 16'b00000_000000_00000;
        tick_overlay[6][11] = 16'b00000_000000_00000;
        tick_overlay[6][12] = 16'b00000_000000_00000;
        tick_overlay[6][13] = 16'b00000_000000_00000;
        tick_overlay[6][14] = 16'b00000_000000_00000;
        tick_overlay[6][15] = 16'b00000_000000_00000;
        tick_overlay[6][16] = 16'b00000_000000_00000;
        tick_overlay[6][17] = 16'b00000_000000_00000;
        tick_overlay[6][18] = 16'b00000_101101_00000;
        tick_overlay[6][19] = 16'b00000_101101_00000;
        tick_overlay[6][20] = 16'b00000_101101_00000;
        tick_overlay[6][21] = 16'b00000_000000_00000;
        tick_overlay[6][22] = 16'b00000_000000_00000;
        tick_overlay[6][23] = 16'b00000_000000_00000;
        tick_overlay[6][24] = 16'b00000_000000_00000;
        tick_overlay[6][25] = 16'b00000_000000_00000;
        tick_overlay[6][26] = 16'b00000_000000_00000;
        tick_overlay[6][27] = 16'b00000_000000_00000;
        tick_overlay[6][28] = 16'b00000_000000_00000;
        tick_overlay[6][29] = 16'b00000_000000_00000;
        tick_overlay[6][30] = 16'b00000_101101_00000;
        tick_overlay[6][31] = 16'b00000_101101_00000;
        tick_overlay[7][0] = 16'b00000_101101_00000;
        tick_overlay[7][1] = 16'b00000_101101_00000;
        tick_overlay[7][2] = 16'b00000_000000_00000;
        tick_overlay[7][3] = 16'b00000_000000_00000;
        tick_overlay[7][4] = 16'b00000_000000_00000;
        tick_overlay[7][5] = 16'b00000_000000_00000;
        tick_overlay[7][6] = 16'b00000_000000_00000;
        tick_overlay[7][7] = 16'b00000_000000_00000;
        tick_overlay[7][8] = 16'b00000_000000_00000;
        tick_overlay[7][9] = 16'b00000_000000_00000;
        tick_overlay[7][10] = 16'b00000_000000_00000;
        tick_overlay[7][11] = 16'b00000_000000_00000;
        tick_overlay[7][12] = 16'b00000_000000_00000;
        tick_overlay[7][13] = 16'b00000_000000_00000;
        tick_overlay[7][14] = 16'b00000_000000_00000;
        tick_overlay[7][15] = 16'b00000_000000_00000;
        tick_overlay[7][16] = 16'b00000_000000_00000;
        tick_overlay[7][17] = 16'b00000_101101_00000;
        tick_overlay[7][18] = 16'b00000_101101_00000;
        tick_overlay[7][19] = 16'b00000_101101_00000;
        tick_overlay[7][20] = 16'b00000_101101_00000;
        tick_overlay[7][21] = 16'b00000_101101_00000;
        tick_overlay[7][22] = 16'b00000_101101_00000;
        tick_overlay[7][23] = 16'b00000_000000_00000;
        tick_overlay[7][24] = 16'b00000_000000_00000;
        tick_overlay[7][25] = 16'b00000_000000_00000;
        tick_overlay[7][26] = 16'b00000_000000_00000;
        tick_overlay[7][27] = 16'b00000_000000_00000;
        tick_overlay[7][28] = 16'b00000_000000_00000;
        tick_overlay[7][29] = 16'b00000_000000_00000;
        tick_overlay[7][30] = 16'b00000_101101_00000;
        tick_overlay[7][31] = 16'b00000_101101_00000;
        tick_overlay[8][0] = 16'b00000_101101_00000;
        tick_overlay[8][1] = 16'b00000_101101_00000;
        tick_overlay[8][2] = 16'b00000_000000_00000;
        tick_overlay[8][3] = 16'b00000_000000_00000;
        tick_overlay[8][4] = 16'b00000_000000_00000;
        tick_overlay[8][5] = 16'b00000_000000_00000;
        tick_overlay[8][6] = 16'b00000_000000_00000;
        tick_overlay[8][7] = 16'b00000_000000_00000;
        tick_overlay[8][8] = 16'b00000_000000_00000;
        tick_overlay[8][9] = 16'b00000_000000_00000;
        tick_overlay[8][10] = 16'b00000_000000_00000;
        tick_overlay[8][11] = 16'b00000_000000_00000;
        tick_overlay[8][12] = 16'b00000_000000_00000;
        tick_overlay[8][13] = 16'b00000_000000_00000;
        tick_overlay[8][14] = 16'b00000_000000_00000;
        tick_overlay[8][15] = 16'b00000_000000_00000;
        tick_overlay[8][16] = 16'b00000_101101_00000;
        tick_overlay[8][17] = 16'b00000_101101_00000;
        tick_overlay[8][18] = 16'b00000_101101_00000;
        tick_overlay[8][19] = 16'b00000_101101_00000;
        tick_overlay[8][20] = 16'b00000_101101_00000;
        tick_overlay[8][21] = 16'b00000_101101_00000;
        tick_overlay[8][22] = 16'b00000_101101_00000;
        tick_overlay[8][23] = 16'b00000_101101_00000;
        tick_overlay[8][24] = 16'b00000_000000_00000;
        tick_overlay[8][25] = 16'b00000_000000_00000;
        tick_overlay[8][26] = 16'b00000_000000_00000;
        tick_overlay[8][27] = 16'b00000_000000_00000;
        tick_overlay[8][28] = 16'b00000_000000_00000;
        tick_overlay[8][29] = 16'b00000_000000_00000;
        tick_overlay[8][30] = 16'b00000_101101_00000;
        tick_overlay[8][31] = 16'b00000_101101_00000;
        tick_overlay[9][0] = 16'b00000_101101_00000;
        tick_overlay[9][1] = 16'b00000_101101_00000;
        tick_overlay[9][2] = 16'b00000_000000_00000;
        tick_overlay[9][3] = 16'b00000_000000_00000;
        tick_overlay[9][4] = 16'b00000_000000_00000;
        tick_overlay[9][5] = 16'b00000_000000_00000;
        tick_overlay[9][6] = 16'b00000_000000_00000;
        tick_overlay[9][7] = 16'b00000_000000_00000;
        tick_overlay[9][8] = 16'b00000_000000_00000;
        tick_overlay[9][9] = 16'b00000_000000_00000;
        tick_overlay[9][10] = 16'b00000_000000_00000;
        tick_overlay[9][11] = 16'b00000_000000_00000;
        tick_overlay[9][12] = 16'b00000_000000_00000;
        tick_overlay[9][13] = 16'b00000_000000_00000;
        tick_overlay[9][14] = 16'b00000_000000_00000;
        tick_overlay[9][15] = 16'b00000_101101_00000;
        tick_overlay[9][16] = 16'b00000_101101_00000;
        tick_overlay[9][17] = 16'b00000_101101_00000;
        tick_overlay[9][18] = 16'b00000_101101_00000;
        tick_overlay[9][19] = 16'b00000_101101_00000;
        tick_overlay[9][20] = 16'b00000_101101_00000;
        tick_overlay[9][21] = 16'b00000_101101_00000;
        tick_overlay[9][22] = 16'b00000_101101_00000;
        tick_overlay[9][23] = 16'b00000_101101_00000;
        tick_overlay[9][24] = 16'b00000_101101_00000;
        tick_overlay[9][25] = 16'b00000_000000_00000;
        tick_overlay[9][26] = 16'b00000_000000_00000;
        tick_overlay[9][27] = 16'b00000_000000_00000;
        tick_overlay[9][28] = 16'b00000_000000_00000;
        tick_overlay[9][29] = 16'b00000_000000_00000;
        tick_overlay[9][30] = 16'b00000_101101_00000;
        tick_overlay[9][31] = 16'b00000_101101_00000;
        tick_overlay[10][0] = 16'b00000_101101_00000;
        tick_overlay[10][1] = 16'b00000_101101_00000;
        tick_overlay[10][2] = 16'b00000_000000_00000;
        tick_overlay[10][3] = 16'b00000_000000_00000;
        tick_overlay[10][4] = 16'b00000_000000_00000;
        tick_overlay[10][5] = 16'b00000_000000_00000;
        tick_overlay[10][6] = 16'b00000_000000_00000;
        tick_overlay[10][7] = 16'b00000_000000_00000;
        tick_overlay[10][8] = 16'b00000_000000_00000;
        tick_overlay[10][9] = 16'b00000_000000_00000;
        tick_overlay[10][10] = 16'b00000_000000_00000;
        tick_overlay[10][11] = 16'b00000_000000_00000;
        tick_overlay[10][12] = 16'b00000_000000_00000;
        tick_overlay[10][13] = 16'b00000_000000_00000;
        tick_overlay[10][14] = 16'b00000_101101_00000;
        tick_overlay[10][15] = 16'b00000_101101_00000;
        tick_overlay[10][16] = 16'b00000_101101_00000;
        tick_overlay[10][17] = 16'b00000_101101_00000;
        tick_overlay[10][18] = 16'b00000_101101_00000;
        tick_overlay[10][19] = 16'b00000_101101_00000;
        tick_overlay[10][20] = 16'b00000_101101_00000;
        tick_overlay[10][21] = 16'b00000_101101_00000;
        tick_overlay[10][22] = 16'b00000_101101_00000;
        tick_overlay[10][23] = 16'b00000_101101_00000;
        tick_overlay[10][24] = 16'b00000_101101_00000;
        tick_overlay[10][25] = 16'b00000_101101_00000;
        tick_overlay[10][26] = 16'b00000_000000_00000;
        tick_overlay[10][27] = 16'b00000_000000_00000;
        tick_overlay[10][28] = 16'b00000_000000_00000;
        tick_overlay[10][29] = 16'b00000_000000_00000;
        tick_overlay[10][30] = 16'b00000_101101_00000;
        tick_overlay[10][31] = 16'b00000_101101_00000;
        tick_overlay[11][0] = 16'b00000_101101_00000;
        tick_overlay[11][1] = 16'b00000_101101_00000;
        tick_overlay[11][2] = 16'b00000_000000_00000;
        tick_overlay[11][3] = 16'b00000_000000_00000;
        tick_overlay[11][4] = 16'b00000_000000_00000;
        tick_overlay[11][5] = 16'b00000_000000_00000;
        tick_overlay[11][6] = 16'b00000_000000_00000;
        tick_overlay[11][7] = 16'b00000_000000_00000;
        tick_overlay[11][8] = 16'b00000_000000_00000;
        tick_overlay[11][9] = 16'b00000_000000_00000;
        tick_overlay[11][10] = 16'b00000_000000_00000;
        tick_overlay[11][11] = 16'b00000_000000_00000;
        tick_overlay[11][12] = 16'b00000_000000_00000;
        tick_overlay[11][13] = 16'b00000_000000_00000;
        tick_overlay[11][14] = 16'b00000_101101_00000;
        tick_overlay[11][15] = 16'b00000_101101_00000;
        tick_overlay[11][16] = 16'b00000_101101_00000;
        tick_overlay[11][17] = 16'b00000_101101_00000;
        tick_overlay[11][18] = 16'b00000_101101_00000;
        tick_overlay[11][19] = 16'b00000_101101_00000;
        tick_overlay[11][20] = 16'b00000_101101_00000;
        tick_overlay[11][21] = 16'b00000_101101_00000;
        tick_overlay[11][22] = 16'b00000_101101_00000;
        tick_overlay[11][23] = 16'b00000_101101_00000;
        tick_overlay[11][24] = 16'b00000_101101_00000;
        tick_overlay[11][25] = 16'b00000_101101_00000;
        tick_overlay[11][26] = 16'b00000_000000_00000;
        tick_overlay[11][27] = 16'b00000_000000_00000;
        tick_overlay[11][28] = 16'b00000_000000_00000;
        tick_overlay[11][29] = 16'b00000_000000_00000;
        tick_overlay[11][30] = 16'b00000_101101_00000;
        tick_overlay[11][31] = 16'b00000_101101_00000;
        tick_overlay[12][0] = 16'b00000_101101_00000;
        tick_overlay[12][1] = 16'b00000_101101_00000;
        tick_overlay[12][2] = 16'b00000_000000_00000;
        tick_overlay[12][3] = 16'b00000_000000_00000;
        tick_overlay[12][4] = 16'b00000_000000_00000;
        tick_overlay[12][5] = 16'b00000_000000_00000;
        tick_overlay[12][6] = 16'b00000_000000_00000;
        tick_overlay[12][7] = 16'b00000_000000_00000;
        tick_overlay[12][8] = 16'b00000_000000_00000;
        tick_overlay[12][9] = 16'b00000_000000_00000;
        tick_overlay[12][10] = 16'b00000_000000_00000;
        tick_overlay[12][11] = 16'b00000_000000_00000;
        tick_overlay[12][12] = 16'b00000_000000_00000;
        tick_overlay[12][13] = 16'b00000_101101_00000;
        tick_overlay[12][14] = 16'b00000_101101_00000;
        tick_overlay[12][15] = 16'b00000_101101_00000;
        tick_overlay[12][16] = 16'b00000_101101_00000;
        tick_overlay[12][17] = 16'b00000_101101_00000;
        tick_overlay[12][18] = 16'b00000_101101_00000;
        tick_overlay[12][19] = 16'b00000_000000_00000;
        tick_overlay[12][20] = 16'b00000_000000_00000;
        tick_overlay[12][21] = 16'b00000_101101_00000;
        tick_overlay[12][22] = 16'b00000_101101_00000;
        tick_overlay[12][23] = 16'b00000_101101_00000;
        tick_overlay[12][24] = 16'b00000_101101_00000;
        tick_overlay[12][25] = 16'b00000_101101_00000;
        tick_overlay[12][26] = 16'b00000_101101_00000;
        tick_overlay[12][27] = 16'b00000_000000_00000;
        tick_overlay[12][28] = 16'b00000_000000_00000;
        tick_overlay[12][29] = 16'b00000_000000_00000;
        tick_overlay[12][30] = 16'b00000_101101_00000;
        tick_overlay[12][31] = 16'b00000_101101_00000;
        tick_overlay[13][0] = 16'b00000_101101_00000;
        tick_overlay[13][1] = 16'b00000_101101_00000;
        tick_overlay[13][2] = 16'b00000_000000_00000;
        tick_overlay[13][3] = 16'b00000_000000_00000;
        tick_overlay[13][4] = 16'b00000_000000_00000;
        tick_overlay[13][5] = 16'b00000_000000_00000;
        tick_overlay[13][6] = 16'b00000_000000_00000;
        tick_overlay[13][7] = 16'b00000_000000_00000;
        tick_overlay[13][8] = 16'b00000_000000_00000;
        tick_overlay[13][9] = 16'b00000_000000_00000;
        tick_overlay[13][10] = 16'b00000_000000_00000;
        tick_overlay[13][11] = 16'b00000_000000_00000;
        tick_overlay[13][12] = 16'b00000_101101_00000;
        tick_overlay[13][13] = 16'b00000_101101_00000;
        tick_overlay[13][14] = 16'b00000_101101_00000;
        tick_overlay[13][15] = 16'b00000_101101_00000;
        tick_overlay[13][16] = 16'b00000_101101_00000;
        tick_overlay[13][17] = 16'b00000_101101_00000;
        tick_overlay[13][18] = 16'b00000_000000_00000;
        tick_overlay[13][19] = 16'b00000_000000_00000;
        tick_overlay[13][20] = 16'b00000_000000_00000;
        tick_overlay[13][21] = 16'b00000_000000_00000;
        tick_overlay[13][22] = 16'b00000_101101_00000;
        tick_overlay[13][23] = 16'b00000_101101_00000;
        tick_overlay[13][24] = 16'b00000_101101_00000;
        tick_overlay[13][25] = 16'b00000_101101_00000;
        tick_overlay[13][26] = 16'b00000_101101_00000;
        tick_overlay[13][27] = 16'b00000_101101_00000;
        tick_overlay[13][28] = 16'b00000_000000_00000;
        tick_overlay[13][29] = 16'b00000_000000_00000;
        tick_overlay[13][30] = 16'b00000_101101_00000;
        tick_overlay[13][31] = 16'b00000_101101_00000;
        tick_overlay[14][0] = 16'b00000_101101_00000;
        tick_overlay[14][1] = 16'b00000_101101_00000;
        tick_overlay[14][2] = 16'b00000_000000_00000;
        tick_overlay[14][3] = 16'b00000_000000_00000;
        tick_overlay[14][4] = 16'b00000_000000_00000;
        tick_overlay[14][5] = 16'b00000_000000_00000;
        tick_overlay[14][6] = 16'b00000_000000_00000;
        tick_overlay[14][7] = 16'b00000_000000_00000;
        tick_overlay[14][8] = 16'b00000_000000_00000;
        tick_overlay[14][9] = 16'b00000_000000_00000;
        tick_overlay[14][10] = 16'b00000_000000_00000;
        tick_overlay[14][11] = 16'b00000_101101_00000;
        tick_overlay[14][12] = 16'b00000_101101_00000;
        tick_overlay[14][13] = 16'b00000_101101_00000;
        tick_overlay[14][14] = 16'b00000_101101_00000;
        tick_overlay[14][15] = 16'b00000_101101_00000;
        tick_overlay[14][16] = 16'b00000_101101_00000;
        tick_overlay[14][17] = 16'b00000_101101_00000;
        tick_overlay[14][18] = 16'b00000_000000_00000;
        tick_overlay[14][19] = 16'b00000_000000_00000;
        tick_overlay[14][20] = 16'b00000_000000_00000;
        tick_overlay[14][21] = 16'b00000_000000_00000;
        tick_overlay[14][22] = 16'b00000_000000_00000;
        tick_overlay[14][23] = 16'b00000_101101_00000;
        tick_overlay[14][24] = 16'b00000_101101_00000;
        tick_overlay[14][25] = 16'b00000_101101_00000;
        tick_overlay[14][26] = 16'b00000_101101_00000;
        tick_overlay[14][27] = 16'b00000_101101_00000;
        tick_overlay[14][28] = 16'b00000_000000_00000;
        tick_overlay[14][29] = 16'b00000_000000_00000;
        tick_overlay[14][30] = 16'b00000_101101_00000;
        tick_overlay[14][31] = 16'b00000_101101_00000;
        tick_overlay[15][0] = 16'b00000_101101_00000;
        tick_overlay[15][1] = 16'b00000_101101_00000;
        tick_overlay[15][2] = 16'b00000_000000_00000;
        tick_overlay[15][3] = 16'b00000_000000_00000;
        tick_overlay[15][4] = 16'b00000_000000_00000;
        tick_overlay[15][5] = 16'b00000_000000_00000;
        tick_overlay[15][6] = 16'b00000_000000_00000;
        tick_overlay[15][7] = 16'b00000_000000_00000;
        tick_overlay[15][8] = 16'b00000_000000_00000;
        tick_overlay[15][9] = 16'b00000_000000_00000;
        tick_overlay[15][10] = 16'b00000_000000_00000;
        tick_overlay[15][11] = 16'b00000_101101_00000;
        tick_overlay[15][12] = 16'b00000_101101_00000;
        tick_overlay[15][13] = 16'b00000_101101_00000;
        tick_overlay[15][14] = 16'b00000_101101_00000;
        tick_overlay[15][15] = 16'b00000_101101_00000;
        tick_overlay[15][16] = 16'b00000_101101_00000;
        tick_overlay[15][17] = 16'b00000_000000_00000;
        tick_overlay[15][18] = 16'b00000_000000_00000;
        tick_overlay[15][19] = 16'b00000_000000_00000;
        tick_overlay[15][20] = 16'b00000_000000_00000;
        tick_overlay[15][21] = 16'b00000_000000_00000;
        tick_overlay[15][22] = 16'b00000_000000_00000;
        tick_overlay[15][23] = 16'b00000_000000_00000;
        tick_overlay[15][24] = 16'b00000_101101_00000;
        tick_overlay[15][25] = 16'b00000_101101_00000;
        tick_overlay[15][26] = 16'b00000_101101_00000;
        tick_overlay[15][27] = 16'b00000_101101_00000;
        tick_overlay[15][28] = 16'b00000_000000_00000;
        tick_overlay[15][29] = 16'b00000_000000_00000;
        tick_overlay[15][30] = 16'b00000_101101_00000;
        tick_overlay[15][31] = 16'b00000_101101_00000;
        tick_overlay[16][0] = 16'b00000_101101_00000;
        tick_overlay[16][1] = 16'b00000_101101_00000;
        tick_overlay[16][2] = 16'b00000_000000_00000;
        tick_overlay[16][3] = 16'b00000_000000_00000;
        tick_overlay[16][4] = 16'b00000_000000_00000;
        tick_overlay[16][5] = 16'b00000_000000_00000;
        tick_overlay[16][6] = 16'b00000_000000_00000;
        tick_overlay[16][7] = 16'b00000_000000_00000;
        tick_overlay[16][8] = 16'b00000_000000_00000;
        tick_overlay[16][9] = 16'b00000_000000_00000;
        tick_overlay[16][10] = 16'b00000_101101_00000;
        tick_overlay[16][11] = 16'b00000_101101_00000;
        tick_overlay[16][12] = 16'b00000_101101_00000;
        tick_overlay[16][13] = 16'b00000_101101_00000;
        tick_overlay[16][14] = 16'b00000_101101_00000;
        tick_overlay[16][15] = 16'b00000_101101_00000;
        tick_overlay[16][16] = 16'b00000_000000_00000;
        tick_overlay[16][17] = 16'b00000_000000_00000;
        tick_overlay[16][18] = 16'b00000_000000_00000;
        tick_overlay[16][19] = 16'b00000_000000_00000;
        tick_overlay[16][20] = 16'b00000_000000_00000;
        tick_overlay[16][21] = 16'b00000_000000_00000;
        tick_overlay[16][22] = 16'b00000_000000_00000;
        tick_overlay[16][23] = 16'b00000_000000_00000;
        tick_overlay[16][24] = 16'b00000_000000_00000;
        tick_overlay[16][25] = 16'b00000_000000_00000;
        tick_overlay[16][26] = 16'b00000_101101_00000;
        tick_overlay[16][27] = 16'b00000_101101_00000;
        tick_overlay[16][28] = 16'b00000_000000_00000;
        tick_overlay[16][29] = 16'b00000_000000_00000;
        tick_overlay[16][30] = 16'b00000_101101_00000;
        tick_overlay[16][31] = 16'b00000_101101_00000;
        tick_overlay[17][0] = 16'b00000_101101_00000;
        tick_overlay[17][1] = 16'b00000_101101_00000;
        tick_overlay[17][2] = 16'b00000_000000_00000;
        tick_overlay[17][3] = 16'b00000_000000_00000;
        tick_overlay[17][4] = 16'b00000_000000_00000;
        tick_overlay[17][5] = 16'b00000_000000_00000;
        tick_overlay[17][6] = 16'b00000_000000_00000;
        tick_overlay[17][7] = 16'b00000_000000_00000;
        tick_overlay[17][8] = 16'b00000_000000_00000;
        tick_overlay[17][9] = 16'b00000_101101_00000;
        tick_overlay[17][10] = 16'b00000_101101_00000;
        tick_overlay[17][11] = 16'b00000_101101_00000;
        tick_overlay[17][12] = 16'b00000_101101_00000;
        tick_overlay[17][13] = 16'b00000_101101_00000;
        tick_overlay[17][14] = 16'b00000_101101_00000;
        tick_overlay[17][15] = 16'b00000_000000_00000;
        tick_overlay[17][16] = 16'b00000_000000_00000;
        tick_overlay[17][17] = 16'b00000_000000_00000;
        tick_overlay[17][18] = 16'b00000_000000_00000;
        tick_overlay[17][19] = 16'b00000_000000_00000;
        tick_overlay[17][20] = 16'b00000_000000_00000;
        tick_overlay[17][21] = 16'b00000_000000_00000;
        tick_overlay[17][22] = 16'b00000_000000_00000;
        tick_overlay[17][23] = 16'b00000_000000_00000;
        tick_overlay[17][24] = 16'b00000_000000_00000;
        tick_overlay[17][25] = 16'b00000_000000_00000;
        tick_overlay[17][26] = 16'b00000_000000_00000;
        tick_overlay[17][27] = 16'b00000_000000_00000;
        tick_overlay[17][28] = 16'b00000_000000_00000;
        tick_overlay[17][29] = 16'b00000_000000_00000;
        tick_overlay[17][30] = 16'b00000_101101_00000;
        tick_overlay[17][31] = 16'b00000_101101_00000;
        tick_overlay[18][0] = 16'b00000_101101_00000;
        tick_overlay[18][1] = 16'b00000_101101_00000;
        tick_overlay[18][2] = 16'b00000_000000_00000;
        tick_overlay[18][3] = 16'b00000_000000_00000;
        tick_overlay[18][4] = 16'b00000_000000_00000;
        tick_overlay[18][5] = 16'b00000_000000_00000;
        tick_overlay[18][6] = 16'b00000_000000_00000;
        tick_overlay[18][7] = 16'b00000_000000_00000;
        tick_overlay[18][8] = 16'b00000_101101_00000;
        tick_overlay[18][9] = 16'b00000_101101_00000;
        tick_overlay[18][10] = 16'b00000_101101_00000;
        tick_overlay[18][11] = 16'b00000_101101_00000;
        tick_overlay[18][12] = 16'b00000_101101_00000;
        tick_overlay[18][13] = 16'b00000_101101_00000;
        tick_overlay[18][14] = 16'b00000_101101_00000;
        tick_overlay[18][15] = 16'b00000_000000_00000;
        tick_overlay[18][16] = 16'b00000_000000_00000;
        tick_overlay[18][17] = 16'b00000_000000_00000;
        tick_overlay[18][18] = 16'b00000_000000_00000;
        tick_overlay[18][19] = 16'b00000_000000_00000;
        tick_overlay[18][20] = 16'b00000_000000_00000;
        tick_overlay[18][21] = 16'b00000_000000_00000;
        tick_overlay[18][22] = 16'b00000_000000_00000;
        tick_overlay[18][23] = 16'b00000_000000_00000;
        tick_overlay[18][24] = 16'b00000_000000_00000;
        tick_overlay[18][25] = 16'b00000_000000_00000;
        tick_overlay[18][26] = 16'b00000_000000_00000;
        tick_overlay[18][27] = 16'b00000_000000_00000;
        tick_overlay[18][28] = 16'b00000_000000_00000;
        tick_overlay[18][29] = 16'b00000_000000_00000;
        tick_overlay[18][30] = 16'b00000_101101_00000;
        tick_overlay[18][31] = 16'b00000_101101_00000;
        tick_overlay[19][0] = 16'b00000_101101_00000;
        tick_overlay[19][1] = 16'b00000_101101_00000;
        tick_overlay[19][2] = 16'b00000_000000_00000;
        tick_overlay[19][3] = 16'b00000_000000_00000;
        tick_overlay[19][4] = 16'b00000_000000_00000;
        tick_overlay[19][5] = 16'b00000_000000_00000;
        tick_overlay[19][6] = 16'b00000_000000_00000;
        tick_overlay[19][7] = 16'b00000_000000_00000;
        tick_overlay[19][8] = 16'b00000_101101_00000;
        tick_overlay[19][9] = 16'b00000_101101_00000;
        tick_overlay[19][10] = 16'b00000_101101_00000;
        tick_overlay[19][11] = 16'b00000_101101_00000;
        tick_overlay[19][12] = 16'b00000_101101_00000;
        tick_overlay[19][13] = 16'b00000_101101_00000;
        tick_overlay[19][14] = 16'b00000_000000_00000;
        tick_overlay[19][15] = 16'b00000_000000_00000;
        tick_overlay[19][16] = 16'b00000_000000_00000;
        tick_overlay[19][17] = 16'b00000_000000_00000;
        tick_overlay[19][18] = 16'b00000_000000_00000;
        tick_overlay[19][19] = 16'b00000_000000_00000;
        tick_overlay[19][20] = 16'b00000_000000_00000;
        tick_overlay[19][21] = 16'b00000_000000_00000;
        tick_overlay[19][22] = 16'b00000_000000_00000;
        tick_overlay[19][23] = 16'b00000_000000_00000;
        tick_overlay[19][24] = 16'b00000_000000_00000;
        tick_overlay[19][25] = 16'b00000_000000_00000;
        tick_overlay[19][26] = 16'b00000_000000_00000;
        tick_overlay[19][27] = 16'b00000_000000_00000;
        tick_overlay[19][28] = 16'b00000_000000_00000;
        tick_overlay[19][29] = 16'b00000_000000_00000;
        tick_overlay[19][30] = 16'b00000_101101_00000;
        tick_overlay[19][31] = 16'b00000_101101_00000;
        tick_overlay[20][0] = 16'b00000_101101_00000;
        tick_overlay[20][1] = 16'b00000_101101_00000;
        tick_overlay[20][2] = 16'b00000_000000_00000;
        tick_overlay[20][3] = 16'b00000_000000_00000;
        tick_overlay[20][4] = 16'b00000_000000_00000;
        tick_overlay[20][5] = 16'b00000_000000_00000;
        tick_overlay[20][6] = 16'b00000_000000_00000;
        tick_overlay[20][7] = 16'b00000_101101_00000;
        tick_overlay[20][8] = 16'b00000_101101_00000;
        tick_overlay[20][9] = 16'b00000_101101_00000;
        tick_overlay[20][10] = 16'b00000_101101_00000;
        tick_overlay[20][11] = 16'b00000_101101_00000;
        tick_overlay[20][12] = 16'b00000_101101_00000;
        tick_overlay[20][13] = 16'b00000_000000_00000;
        tick_overlay[20][14] = 16'b00000_000000_00000;
        tick_overlay[20][15] = 16'b00000_000000_00000;
        tick_overlay[20][16] = 16'b00000_000000_00000;
        tick_overlay[20][17] = 16'b00000_000000_00000;
        tick_overlay[20][18] = 16'b00000_000000_00000;
        tick_overlay[20][19] = 16'b00000_000000_00000;
        tick_overlay[20][20] = 16'b00000_000000_00000;
        tick_overlay[20][21] = 16'b00000_000000_00000;
        tick_overlay[20][22] = 16'b00000_000000_00000;
        tick_overlay[20][23] = 16'b00000_000000_00000;
        tick_overlay[20][24] = 16'b00000_000000_00000;
        tick_overlay[20][25] = 16'b00000_000000_00000;
        tick_overlay[20][26] = 16'b00000_000000_00000;
        tick_overlay[20][27] = 16'b00000_000000_00000;
        tick_overlay[20][28] = 16'b00000_000000_00000;
        tick_overlay[20][29] = 16'b00000_000000_00000;
        tick_overlay[20][30] = 16'b00000_101101_00000;
        tick_overlay[20][31] = 16'b00000_101101_00000;
        tick_overlay[21][0] = 16'b00000_101101_00000;
        tick_overlay[21][1] = 16'b00000_101101_00000;
        tick_overlay[21][2] = 16'b00000_000000_00000;
        tick_overlay[21][3] = 16'b00000_000000_00000;
        tick_overlay[21][4] = 16'b00000_000000_00000;
        tick_overlay[21][5] = 16'b00000_000000_00000;
        tick_overlay[21][6] = 16'b00000_101101_00000;
        tick_overlay[21][7] = 16'b00000_101101_00000;
        tick_overlay[21][8] = 16'b00000_101101_00000;
        tick_overlay[21][9] = 16'b00000_101101_00000;
        tick_overlay[21][10] = 16'b00000_101101_00000;
        tick_overlay[21][11] = 16'b00000_101101_00000;
        tick_overlay[21][12] = 16'b00000_000000_00000;
        tick_overlay[21][13] = 16'b00000_000000_00000;
        tick_overlay[21][14] = 16'b00000_000000_00000;
        tick_overlay[21][15] = 16'b00000_000000_00000;
        tick_overlay[21][16] = 16'b00000_000000_00000;
        tick_overlay[21][17] = 16'b00000_000000_00000;
        tick_overlay[21][18] = 16'b00000_000000_00000;
        tick_overlay[21][19] = 16'b00000_000000_00000;
        tick_overlay[21][20] = 16'b00000_000000_00000;
        tick_overlay[21][21] = 16'b00000_000000_00000;
        tick_overlay[21][22] = 16'b00000_000000_00000;
        tick_overlay[21][23] = 16'b00000_000000_00000;
        tick_overlay[21][24] = 16'b00000_000000_00000;
        tick_overlay[21][25] = 16'b00000_000000_00000;
        tick_overlay[21][26] = 16'b00000_000000_00000;
        tick_overlay[21][27] = 16'b00000_000000_00000;
        tick_overlay[21][28] = 16'b00000_000000_00000;
        tick_overlay[21][29] = 16'b00000_000000_00000;
        tick_overlay[21][30] = 16'b00000_101101_00000;
        tick_overlay[21][31] = 16'b00000_101101_00000;
        tick_overlay[22][0] = 16'b00000_101101_00000;
        tick_overlay[22][1] = 16'b00000_101101_00000;
        tick_overlay[22][2] = 16'b00000_000000_00000;
        tick_overlay[22][3] = 16'b00000_000000_00000;
        tick_overlay[22][4] = 16'b00000_000000_00000;
        tick_overlay[22][5] = 16'b00000_101101_00000;
        tick_overlay[22][6] = 16'b00000_101101_00000;
        tick_overlay[22][7] = 16'b00000_101101_00000;
        tick_overlay[22][8] = 16'b00000_101101_00000;
        tick_overlay[22][9] = 16'b00000_101101_00000;
        tick_overlay[22][10] = 16'b00000_101101_00000;
        tick_overlay[22][11] = 16'b00000_000000_00000;
        tick_overlay[22][12] = 16'b00000_000000_00000;
        tick_overlay[22][13] = 16'b00000_000000_00000;
        tick_overlay[22][14] = 16'b00000_000000_00000;
        tick_overlay[22][15] = 16'b00000_000000_00000;
        tick_overlay[22][16] = 16'b00000_000000_00000;
        tick_overlay[22][17] = 16'b00000_000000_00000;
        tick_overlay[22][18] = 16'b00000_000000_00000;
        tick_overlay[22][19] = 16'b00000_000000_00000;
        tick_overlay[22][20] = 16'b00000_000000_00000;
        tick_overlay[22][21] = 16'b00000_000000_00000;
        tick_overlay[22][22] = 16'b00000_000000_00000;
        tick_overlay[22][23] = 16'b00000_000000_00000;
        tick_overlay[22][24] = 16'b00000_000000_00000;
        tick_overlay[22][25] = 16'b00000_000000_00000;
        tick_overlay[22][26] = 16'b00000_000000_00000;
        tick_overlay[22][27] = 16'b00000_000000_00000;
        tick_overlay[22][28] = 16'b00000_000000_00000;
        tick_overlay[22][29] = 16'b00000_000000_00000;
        tick_overlay[22][30] = 16'b00000_101101_00000;
        tick_overlay[22][31] = 16'b00000_101101_00000;
        tick_overlay[23][0] = 16'b00000_101101_00000;
        tick_overlay[23][1] = 16'b00000_101101_00000;
        tick_overlay[23][2] = 16'b00000_000000_00000;
        tick_overlay[23][3] = 16'b00000_000000_00000;
        tick_overlay[23][4] = 16'b00000_000000_00000;
        tick_overlay[23][5] = 16'b00000_101101_00000;
        tick_overlay[23][6] = 16'b00000_101101_00000;
        tick_overlay[23][7] = 16'b00000_101101_00000;
        tick_overlay[23][8] = 16'b00000_101101_00000;
        tick_overlay[23][9] = 16'b00000_101101_00000;
        tick_overlay[23][10] = 16'b00000_000000_00000;
        tick_overlay[23][11] = 16'b00000_000000_00000;
        tick_overlay[23][12] = 16'b00000_000000_00000;
        tick_overlay[23][13] = 16'b00000_000000_00000;
        tick_overlay[23][14] = 16'b00000_000000_00000;
        tick_overlay[23][15] = 16'b00000_000000_00000;
        tick_overlay[23][16] = 16'b00000_000000_00000;
        tick_overlay[23][17] = 16'b00000_000000_00000;
        tick_overlay[23][18] = 16'b00000_000000_00000;
        tick_overlay[23][19] = 16'b00000_000000_00000;
        tick_overlay[23][20] = 16'b00000_000000_00000;
        tick_overlay[23][21] = 16'b00000_000000_00000;
        tick_overlay[23][22] = 16'b00000_000000_00000;
        tick_overlay[23][23] = 16'b00000_000000_00000;
        tick_overlay[23][24] = 16'b00000_000000_00000;
        tick_overlay[23][25] = 16'b00000_000000_00000;
        tick_overlay[23][26] = 16'b00000_000000_00000;
        tick_overlay[23][27] = 16'b00000_000000_00000;
        tick_overlay[23][28] = 16'b00000_000000_00000;
        tick_overlay[23][29] = 16'b00000_000000_00000;
        tick_overlay[23][30] = 16'b00000_101101_00000;
        tick_overlay[23][31] = 16'b00000_101101_00000;
        tick_overlay[24][0] = 16'b00000_101101_00000;
        tick_overlay[24][1] = 16'b00000_101101_00000;
        tick_overlay[24][2] = 16'b00000_000000_00000;
        tick_overlay[24][3] = 16'b00000_000000_00000;
        tick_overlay[24][4] = 16'b00000_101101_00000;
        tick_overlay[24][5] = 16'b00000_101101_00000;
        tick_overlay[24][6] = 16'b00000_101101_00000;
        tick_overlay[24][7] = 16'b00000_101101_00000;
        tick_overlay[24][8] = 16'b00000_101101_00000;
        tick_overlay[24][9] = 16'b00000_000000_00000;
        tick_overlay[24][10] = 16'b00000_000000_00000;
        tick_overlay[24][11] = 16'b00000_000000_00000;
        tick_overlay[24][12] = 16'b00000_000000_00000;
        tick_overlay[24][13] = 16'b00000_000000_00000;
        tick_overlay[24][14] = 16'b00000_000000_00000;
        tick_overlay[24][15] = 16'b00000_000000_00000;
        tick_overlay[24][16] = 16'b00000_000000_00000;
        tick_overlay[24][17] = 16'b00000_000000_00000;
        tick_overlay[24][18] = 16'b00000_000000_00000;
        tick_overlay[24][19] = 16'b00000_000000_00000;
        tick_overlay[24][20] = 16'b00000_000000_00000;
        tick_overlay[24][21] = 16'b00000_000000_00000;
        tick_overlay[24][22] = 16'b00000_000000_00000;
        tick_overlay[24][23] = 16'b00000_000000_00000;
        tick_overlay[24][24] = 16'b00000_000000_00000;
        tick_overlay[24][25] = 16'b00000_000000_00000;
        tick_overlay[24][26] = 16'b00000_000000_00000;
        tick_overlay[24][27] = 16'b00000_000000_00000;
        tick_overlay[24][28] = 16'b00000_000000_00000;
        tick_overlay[24][29] = 16'b00000_000000_00000;
        tick_overlay[24][30] = 16'b00000_101101_00000;
        tick_overlay[24][31] = 16'b00000_101101_00000;
        tick_overlay[25][0] = 16'b00000_101101_00000;
        tick_overlay[25][1] = 16'b00000_101101_00000;
        tick_overlay[25][2] = 16'b00000_000000_00000;
        tick_overlay[25][3] = 16'b00000_000000_00000;
        tick_overlay[25][4] = 16'b00000_101101_00000;
        tick_overlay[25][5] = 16'b00000_101101_00000;
        tick_overlay[25][6] = 16'b00000_101101_00000;
        tick_overlay[25][7] = 16'b00000_101101_00000;
        tick_overlay[25][8] = 16'b00000_000000_00000;
        tick_overlay[25][9] = 16'b00000_000000_00000;
        tick_overlay[25][10] = 16'b00000_000000_00000;
        tick_overlay[25][11] = 16'b00000_000000_00000;
        tick_overlay[25][12] = 16'b00000_000000_00000;
        tick_overlay[25][13] = 16'b00000_000000_00000;
        tick_overlay[25][14] = 16'b00000_000000_00000;
        tick_overlay[25][15] = 16'b00000_000000_00000;
        tick_overlay[25][16] = 16'b00000_000000_00000;
        tick_overlay[25][17] = 16'b00000_000000_00000;
        tick_overlay[25][18] = 16'b00000_000000_00000;
        tick_overlay[25][19] = 16'b00000_000000_00000;
        tick_overlay[25][20] = 16'b00000_000000_00000;
        tick_overlay[25][21] = 16'b00000_000000_00000;
        tick_overlay[25][22] = 16'b00000_000000_00000;
        tick_overlay[25][23] = 16'b00000_000000_00000;
        tick_overlay[25][24] = 16'b00000_000000_00000;
        tick_overlay[25][25] = 16'b00000_000000_00000;
        tick_overlay[25][26] = 16'b00000_000000_00000;
        tick_overlay[25][27] = 16'b00000_000000_00000;
        tick_overlay[25][28] = 16'b00000_000000_00000;
        tick_overlay[25][29] = 16'b00000_000000_00000;
        tick_overlay[25][30] = 16'b00000_101101_00000;
        tick_overlay[25][31] = 16'b00000_101101_00000;
        tick_overlay[26][0] = 16'b00000_101101_00000;
        tick_overlay[26][1] = 16'b00000_101101_00000;
        tick_overlay[26][2] = 16'b00000_000000_00000;
        tick_overlay[26][3] = 16'b00000_000000_00000;
        tick_overlay[26][4] = 16'b00000_101101_00000;
        tick_overlay[26][5] = 16'b00000_101101_00000;
        tick_overlay[26][6] = 16'b00000_101101_00000;
        tick_overlay[26][7] = 16'b00000_000000_00000;
        tick_overlay[26][8] = 16'b00000_000000_00000;
        tick_overlay[26][9] = 16'b00000_000000_00000;
        tick_overlay[26][10] = 16'b00000_000000_00000;
        tick_overlay[26][11] = 16'b00000_000000_00000;
        tick_overlay[26][12] = 16'b00000_000000_00000;
        tick_overlay[26][13] = 16'b00000_000000_00000;
        tick_overlay[26][14] = 16'b00000_000000_00000;
        tick_overlay[26][15] = 16'b00000_000000_00000;
        tick_overlay[26][16] = 16'b00000_000000_00000;
        tick_overlay[26][17] = 16'b00000_000000_00000;
        tick_overlay[26][18] = 16'b00000_000000_00000;
        tick_overlay[26][19] = 16'b00000_000000_00000;
        tick_overlay[26][20] = 16'b00000_000000_00000;
        tick_overlay[26][21] = 16'b00000_000000_00000;
        tick_overlay[26][22] = 16'b00000_000000_00000;
        tick_overlay[26][23] = 16'b00000_000000_00000;
        tick_overlay[26][24] = 16'b00000_000000_00000;
        tick_overlay[26][25] = 16'b00000_000000_00000;
        tick_overlay[26][26] = 16'b00000_000000_00000;
        tick_overlay[26][27] = 16'b00000_000000_00000;
        tick_overlay[26][28] = 16'b00000_000000_00000;
        tick_overlay[26][29] = 16'b00000_000000_00000;
        tick_overlay[26][30] = 16'b00000_101101_00000;
        tick_overlay[26][31] = 16'b00000_101101_00000;
        tick_overlay[27][0] = 16'b00000_101101_00000;
        tick_overlay[27][1] = 16'b00000_101101_00000;
        tick_overlay[27][2] = 16'b00000_000000_00000;
        tick_overlay[27][3] = 16'b00000_000000_00000;
        tick_overlay[27][4] = 16'b00000_101101_00000;
        tick_overlay[27][5] = 16'b00000_101101_00000;
        tick_overlay[27][6] = 16'b00000_000000_00000;
        tick_overlay[27][7] = 16'b00000_000000_00000;
        tick_overlay[27][8] = 16'b00000_000000_00000;
        tick_overlay[27][9] = 16'b00000_000000_00000;
        tick_overlay[27][10] = 16'b00000_000000_00000;
        tick_overlay[27][11] = 16'b00000_000000_00000;
        tick_overlay[27][12] = 16'b00000_000000_00000;
        tick_overlay[27][13] = 16'b00000_000000_00000;
        tick_overlay[27][14] = 16'b00000_000000_00000;
        tick_overlay[27][15] = 16'b00000_000000_00000;
        tick_overlay[27][16] = 16'b00000_000000_00000;
        tick_overlay[27][17] = 16'b00000_000000_00000;
        tick_overlay[27][18] = 16'b00000_000000_00000;
        tick_overlay[27][19] = 16'b00000_000000_00000;
        tick_overlay[27][20] = 16'b00000_000000_00000;
        tick_overlay[27][21] = 16'b00000_000000_00000;
        tick_overlay[27][22] = 16'b00000_000000_00000;
        tick_overlay[27][23] = 16'b00000_000000_00000;
        tick_overlay[27][24] = 16'b00000_000000_00000;
        tick_overlay[27][25] = 16'b00000_000000_00000;
        tick_overlay[27][26] = 16'b00000_000000_00000;
        tick_overlay[27][27] = 16'b00000_000000_00000;
        tick_overlay[27][28] = 16'b00000_000000_00000;
        tick_overlay[27][29] = 16'b00000_000000_00000;
        tick_overlay[27][30] = 16'b00000_101101_00000;
        tick_overlay[27][31] = 16'b00000_101101_00000;
        tick_overlay[28][0] = 16'b00000_101101_00000;
        tick_overlay[28][1] = 16'b00000_101101_00000;
        tick_overlay[28][2] = 16'b00000_000000_00000;
        tick_overlay[28][3] = 16'b00000_000000_00000;
        tick_overlay[28][4] = 16'b00000_000000_00000;
        tick_overlay[28][5] = 16'b00000_000000_00000;
        tick_overlay[28][6] = 16'b00000_000000_00000;
        tick_overlay[28][7] = 16'b00000_000000_00000;
        tick_overlay[28][8] = 16'b00000_000000_00000;
        tick_overlay[28][9] = 16'b00000_000000_00000;
        tick_overlay[28][10] = 16'b00000_000000_00000;
        tick_overlay[28][11] = 16'b00000_000000_00000;
        tick_overlay[28][12] = 16'b00000_000000_00000;
        tick_overlay[28][13] = 16'b00000_000000_00000;
        tick_overlay[28][14] = 16'b00000_000000_00000;
        tick_overlay[28][15] = 16'b00000_000000_00000;
        tick_overlay[28][16] = 16'b00000_000000_00000;
        tick_overlay[28][17] = 16'b00000_000000_00000;
        tick_overlay[28][18] = 16'b00000_000000_00000;
        tick_overlay[28][19] = 16'b00000_000000_00000;
        tick_overlay[28][20] = 16'b00000_000000_00000;
        tick_overlay[28][21] = 16'b00000_000000_00000;
        tick_overlay[28][22] = 16'b00000_000000_00000;
        tick_overlay[28][23] = 16'b00000_000000_00000;
        tick_overlay[28][24] = 16'b00000_000000_00000;
        tick_overlay[28][25] = 16'b00000_000000_00000;
        tick_overlay[28][26] = 16'b00000_000000_00000;
        tick_overlay[28][27] = 16'b00000_000000_00000;
        tick_overlay[28][28] = 16'b00000_000000_00000;
        tick_overlay[28][29] = 16'b00000_000000_00000;
        tick_overlay[28][30] = 16'b00000_101101_00000;
        tick_overlay[28][31] = 16'b00000_101101_00000;
        tick_overlay[29][0] = 16'b00000_101101_00000;
        tick_overlay[29][1] = 16'b00000_101101_00000;
        tick_overlay[29][2] = 16'b00000_000000_00000;
        tick_overlay[29][3] = 16'b00000_000000_00000;
        tick_overlay[29][4] = 16'b00000_000000_00000;
        tick_overlay[29][5] = 16'b00000_000000_00000;
        tick_overlay[29][6] = 16'b00000_000000_00000;
        tick_overlay[29][7] = 16'b00000_000000_00000;
        tick_overlay[29][8] = 16'b00000_000000_00000;
        tick_overlay[29][9] = 16'b00000_000000_00000;
        tick_overlay[29][10] = 16'b00000_000000_00000;
        tick_overlay[29][11] = 16'b00000_000000_00000;
        tick_overlay[29][12] = 16'b00000_000000_00000;
        tick_overlay[29][13] = 16'b00000_000000_00000;
        tick_overlay[29][14] = 16'b00000_000000_00000;
        tick_overlay[29][15] = 16'b00000_000000_00000;
        tick_overlay[29][16] = 16'b00000_000000_00000;
        tick_overlay[29][17] = 16'b00000_000000_00000;
        tick_overlay[29][18] = 16'b00000_000000_00000;
        tick_overlay[29][19] = 16'b00000_000000_00000;
        tick_overlay[29][20] = 16'b00000_000000_00000;
        tick_overlay[29][21] = 16'b00000_000000_00000;
        tick_overlay[29][22] = 16'b00000_000000_00000;
        tick_overlay[29][23] = 16'b00000_000000_00000;
        tick_overlay[29][24] = 16'b00000_000000_00000;
        tick_overlay[29][25] = 16'b00000_000000_00000;
        tick_overlay[29][26] = 16'b00000_000000_00000;
        tick_overlay[29][27] = 16'b00000_000000_00000;
        tick_overlay[29][28] = 16'b00000_000000_00000;
        tick_overlay[29][29] = 16'b00000_000000_00000;
        tick_overlay[29][30] = 16'b00000_101101_00000;
        tick_overlay[29][31] = 16'b00000_101101_00000;
        tick_overlay[30][0] = 16'b00000_101101_00000;
        tick_overlay[30][1] = 16'b00000_101101_00000;
        tick_overlay[30][2] = 16'b00000_101101_00000;
        tick_overlay[30][3] = 16'b00000_101101_00000;
        tick_overlay[30][4] = 16'b00000_101101_00000;
        tick_overlay[30][5] = 16'b00000_101101_00000;
        tick_overlay[30][6] = 16'b00000_101101_00000;
        tick_overlay[30][7] = 16'b00000_101101_00000;
        tick_overlay[30][8] = 16'b00000_101101_00000;
        tick_overlay[30][9] = 16'b00000_101101_00000;
        tick_overlay[30][10] = 16'b00000_101101_00000;
        tick_overlay[30][11] = 16'b00000_101101_00000;
        tick_overlay[30][12] = 16'b00000_101101_00000;
        tick_overlay[30][13] = 16'b00000_101101_00000;
        tick_overlay[30][14] = 16'b00000_101101_00000;
        tick_overlay[30][15] = 16'b00000_101101_00000;
        tick_overlay[30][16] = 16'b00000_101101_00000;
        tick_overlay[30][17] = 16'b00000_101101_00000;
        tick_overlay[30][18] = 16'b00000_101101_00000;
        tick_overlay[30][19] = 16'b00000_101101_00000;
        tick_overlay[30][20] = 16'b00000_101101_00000;
        tick_overlay[30][21] = 16'b00000_101101_00000;
        tick_overlay[30][22] = 16'b00000_101101_00000;
        tick_overlay[30][23] = 16'b00000_101101_00000;
        tick_overlay[30][24] = 16'b00000_101101_00000;
        tick_overlay[30][25] = 16'b00000_101101_00000;
        tick_overlay[30][26] = 16'b00000_101101_00000;
        tick_overlay[30][27] = 16'b00000_101101_00000;
        tick_overlay[30][28] = 16'b00000_101101_00000;
        tick_overlay[30][29] = 16'b00000_101101_00000;
        tick_overlay[30][30] = 16'b00000_101101_00000;
        tick_overlay[30][31] = 16'b00000_101101_00000;
        tick_overlay[31][0] = 16'b00000_101101_00000;
        tick_overlay[31][1] = 16'b00000_101101_00000;
        tick_overlay[31][2] = 16'b00000_101101_00000;
        tick_overlay[31][3] = 16'b00000_101101_00000;
        tick_overlay[31][4] = 16'b00000_101101_00000;
        tick_overlay[31][5] = 16'b00000_101101_00000;
        tick_overlay[31][6] = 16'b00000_101101_00000;
        tick_overlay[31][7] = 16'b00000_101101_00000;
        tick_overlay[31][8] = 16'b00000_101101_00000;
        tick_overlay[31][9] = 16'b00000_101101_00000;
        tick_overlay[31][10] = 16'b00000_101101_00000;
        tick_overlay[31][11] = 16'b00000_101101_00000;
        tick_overlay[31][12] = 16'b00000_101101_00000;
        tick_overlay[31][13] = 16'b00000_101101_00000;
        tick_overlay[31][14] = 16'b00000_101101_00000;
        tick_overlay[31][15] = 16'b00000_101101_00000;
        tick_overlay[31][16] = 16'b00000_101101_00000;
        tick_overlay[31][17] = 16'b00000_101101_00000;
        tick_overlay[31][18] = 16'b00000_101101_00000;
        tick_overlay[31][19] = 16'b00000_101101_00000;
        tick_overlay[31][20] = 16'b00000_101101_00000;
        tick_overlay[31][21] = 16'b00000_101101_00000;
        tick_overlay[31][22] = 16'b00000_101101_00000;
        tick_overlay[31][23] = 16'b00000_101101_00000;
        tick_overlay[31][24] = 16'b00000_101101_00000;
        tick_overlay[31][25] = 16'b00000_101101_00000;
        tick_overlay[31][26] = 16'b00000_101101_00000;
        tick_overlay[31][27] = 16'b00000_101101_00000;
        tick_overlay[31][28] = 16'b00000_101101_00000;
        tick_overlay[31][29] = 16'b00000_101101_00000;
        tick_overlay[31][30] = 16'b00000_101101_00000;
        tick_overlay[31][31] = 16'b00000_101101_00000;


end



always @(posedge clk) begin

    if (rot_x >= item_1_x_offset && rot_x < item_1_x_offset+32 &&
        rot_y >= item_1_y_offset && rot_y < item_1_y_offset+32) begin
        
        case (item_1_id)
        2'b00: begin
            oled_data <= !orders_done[2] ? (chicken_rice[31 - (rot_y - item_1_y_offset)][31 - (rot_x - item_1_x_offset)]) : ( (chicken_rice_dim[31 - (rot_y - item_1_y_offset)][31 - (rot_x - item_1_x_offset)]) | tick_overlay[31 - (rot_y - item_1_y_offset)][31 - (rot_x - item_1_x_offset)]);
        end
        2'b01: begin
            oled_data <= !orders_done[2] ? (onion_soup[31 - (rot_y - item_1_y_offset)][31 - (rot_x - item_1_x_offset)]) : ( (onion_soup_dim[31 - (rot_y - item_1_y_offset)][31 - (rot_x - item_1_x_offset)]) | tick_overlay[31 - (rot_y - item_1_y_offset)][31 - (rot_x - item_1_x_offset)]);
        end
        2'b10: begin
            oled_data <= !orders_done[2] ? (tomato_soup[31 - (rot_y - item_1_y_offset)][31 - (rot_x - item_1_x_offset)]) : ( (tomato_soup_dim[31 - (rot_y - item_1_y_offset)][31 - (rot_x - item_1_x_offset)]) | tick_overlay[31 - (rot_y - item_1_y_offset)][31 - (rot_x - item_1_x_offset)]);
        end
        2'b11: begin
            oled_data <= !orders_done[2] ? (tomato_rice[31 - (rot_y - item_1_y_offset)][31 - (rot_x - item_1_x_offset)]) : ( (tomato_rice_dim[31 - (rot_y - item_1_y_offset)][31 - (rot_x - item_1_x_offset)]) | tick_overlay[31 - (rot_y - item_1_y_offset)][31 - (rot_x - item_1_x_offset)]);
        end
        endcase
    end


    else if (rot_x >= item_2_x_offset && rot_x < item_2_x_offset+32 && rot_y >= item_2_y_offset && rot_y < item_2_y_offset+32) begin
        case (item_2_id)
        2'b00: begin
            oled_data <= !orders_done[1] ? (chicken_rice[31 - (rot_y - item_2_y_offset)][31 - (rot_x - item_2_x_offset)]) : ( (chicken_rice_dim[31 - (rot_y - item_2_y_offset)][31 - (rot_x - item_2_x_offset)]) | tick_overlay[31 - (rot_y - item_2_y_offset)][31 - (rot_x - item_2_x_offset)]);
        end
        2'b01: begin
            oled_data <= !orders_done[1] ? (onion_soup[31 - (rot_y - item_2_y_offset)][31 - (rot_x - item_2_x_offset)]) : ( (onion_soup_dim[31 - (rot_y - item_2_y_offset)][31 - (rot_x - item_2_x_offset)]) | tick_overlay[31 - (rot_y - item_2_y_offset)][31 - (rot_x - item_2_x_offset)]);
        end
        2'b10: begin
            oled_data <= !orders_done[1] ? (tomato_soup[31 - (rot_y - item_2_y_offset)][31 - (rot_x - item_2_x_offset)]) : ( (tomato_soup_dim[31 - (rot_y - item_2_y_offset)][31 - (rot_x - item_2_x_offset)]) | tick_overlay[31 - (rot_y - item_2_y_offset)][31 - (rot_x - item_2_x_offset)]);
        end
        2'b11: begin
            oled_data <= !orders_done[1] ? (tomato_rice[31 - (rot_y - item_2_y_offset)][31 - (rot_x - item_2_x_offset)]) : ( (tomato_rice_dim[31 - (rot_y - item_2_y_offset)][31 - (rot_x - item_2_x_offset)]) | tick_overlay[31 - (rot_y - item_2_y_offset)][31 - (rot_x - item_2_x_offset)]);
        end
        endcase
    end


    else if (rot_x >= item_3_x_offset && rot_x < item_3_x_offset+32 && rot_y >= item_3_y_offset && rot_y < item_3_y_offset+32) begin
        case (item_3_id)
        2'b00: begin
            oled_data <= !orders_done[0] ? (chicken_rice[31 - (rot_y - item_3_y_offset)][31 - (rot_x - item_3_x_offset)]) : ( (chicken_rice_dim[31 - (rot_y - item_3_y_offset)][31 - (rot_x - item_3_x_offset)]) | tick_overlay[31 - (rot_y - item_3_y_offset)][31 - (rot_x - item_3_x_offset)]);
        end
        2'b01: begin
            oled_data <= !orders_done[0] ? (onion_soup[31 - (rot_y - item_3_y_offset)][31 - (rot_x - item_3_x_offset)]) : ( (onion_soup_dim[31 - (rot_y - item_3_y_offset)][31 - (rot_x - item_3_x_offset)]) | tick_overlay[31 - (rot_y - item_3_y_offset)][31 - (rot_x - item_3_x_offset)]);
        end
        2'b10: begin
            oled_data <= !orders_done[0] ? (tomato_soup[31 - (rot_y - item_3_y_offset)][31 - (rot_x - item_3_x_offset)]) : ( (tomato_soup_dim[31 - (rot_y - item_3_y_offset)][31 - (rot_x - item_3_x_offset)]) | tick_overlay[31 - (rot_y - item_3_y_offset)][31 - (rot_x - item_3_x_offset)]);
        end
        2'b11: begin
            oled_data <= !orders_done[0] ? (tomato_rice[31 - (rot_y - item_3_y_offset)][31 - (rot_x - item_3_x_offset)]) : ( (tomato_rice_dim[31 - (rot_y - item_3_y_offset)][31 - (rot_x - item_3_x_offset)]) | tick_overlay[31 - (rot_y - item_3_y_offset)][31 - (rot_x - item_3_x_offset)]);
        end
        endcase
    end


    else if (rot_x >= ingredient_text_x_offset && rot_x < ingredient_text_x_offset+80 && rot_y >= ingredient_text_y_offset && rot_y < ingredient_text_y_offset+17) begin
        oled_data <= ingredient_text[16 - (rot_y - ingredient_text_y_offset)][79 - (rot_x - ingredient_text_x_offset)];
    end

    else if (rot_x >= holding_ingredient_x_offset && rot_x < holding_ingredient_x_offset+15 && rot_y >= holding_ingredient_y_offset && rot_y < holding_ingredient_y_offset+15) begin
        case (holding_ingredient_id)
            12'b000_000_000_000: oled_data <= 0;
            12'b000_000_000_001: oled_data <= onion_boiled[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b000_000_000_010: oled_data <= onion_chopped[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b000_000_000_100: oled_data <= onion_raw[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b000_000_000_011: oled_data <= onion_boiled_chopped [14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b000_000_001_000: oled_data <= rice_boiled[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b000_000_010_000: oled_data <= rice_chopped[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b000_000_100_000: oled_data <= rice_raw[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b000_000_011_000: oled_data <= rice_boiled_chopped[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b000_001_000_000: oled_data <= tomato_boiled[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b000_010_000_000: oled_data <= tomato_chopped[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b000_100_000_000: oled_data <= tomato_raw[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b000_011_000_000: oled_data <= tomato_boiled_chopped[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b001_000_000_000: oled_data <= chicken_boiled[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b010_000_000_000: oled_data <= chicken_chopped[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b100_000_000_000: oled_data <= chicken_raw[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            12'b011_000_000_000: oled_data <= chicken_boiled_chopped[14-(rot_y-holding_ingredient_y_offset)][14-(rot_x-holding_ingredient_x_offset)];
            default: oled_data <= 0;
        endcase
    end

    else if (rot_x >= item_1_ingredient_1_x_offset && rot_x < item_1_ingredient_1_x_offset+15 && rot_y >= item_1_ingredient_1_y_offset && rot_y < item_1_ingredient_1_y_offset+15) begin
        case (item_1_id)
            2'b00: oled_data <= chicken_boiled_chopped[14-(rot_y-item_1_ingredient_1_y_offset)][14-(rot_x-item_1_ingredient_1_x_offset)];
            2'b01: oled_data <= onion_boiled[14-(rot_y-item_1_ingredient_1_y_offset)][14-(rot_x-item_1_ingredient_1_x_offset)];
            2'b10: oled_data <= tomato_boiled[14-(rot_y-item_1_ingredient_1_y_offset)][14-(rot_x-item_1_ingredient_1_x_offset)];
            2'b11: oled_data <= tomato_boiled[14-(rot_y-item_1_ingredient_1_y_offset)][14-(rot_x-item_1_ingredient_1_x_offset)];
        endcase
    end


    else if (rot_x >= item_1_ingredient_2_x_offset && rot_x < item_1_ingredient_2_x_offset+15 && rot_y >= item_1_ingredient_2_y_offset && rot_y < item_1_ingredient_2_y_offset+15) begin
        case (item_1_id)
            2'b00: oled_data <= rice_boiled[14-(rot_y-item_1_ingredient_2_y_offset)][14-(rot_x-item_1_ingredient_2_x_offset)];
            2'b01: oled_data <= cross[14-(rot_y-item_1_ingredient_2_y_offset)][14-(rot_x-item_1_ingredient_2_x_offset)];
            2'b10: oled_data <= cross[14-(rot_y-item_1_ingredient_2_y_offset)][14-(rot_x-item_1_ingredient_2_x_offset)];
            2'b11: oled_data <= rice_boiled[14-(rot_y-item_1_ingredient_2_y_offset)][14-(rot_x-item_1_ingredient_2_x_offset)];
        endcase
    end


    else if (rot_x >= item_2_ingredient_1_x_offset && rot_x < item_2_ingredient_1_x_offset+15 && rot_y >= item_2_ingredient_1_y_offset && rot_y < item_2_ingredient_1_y_offset+15) begin
        case (item_2_id)
            2'b00: oled_data <= chicken_boiled_chopped[14-(rot_y-item_2_ingredient_1_y_offset)][14-(rot_x-item_2_ingredient_1_x_offset)];
            2'b01: oled_data <= onion_boiled[14-(rot_y-item_2_ingredient_1_y_offset)][14-(rot_x-item_2_ingredient_1_x_offset)];
            2'b10: oled_data <= tomato_boiled[14-(rot_y-item_2_ingredient_1_y_offset)][14-(rot_x-item_2_ingredient_1_x_offset)];
            2'b11: oled_data <= tomato_boiled[14-(rot_y-item_2_ingredient_1_y_offset)][14-(rot_x-item_2_ingredient_1_x_offset)];
        endcase
    end

    else if (rot_x >= item_2_ingredient_2_x_offset && rot_x < item_2_ingredient_2_x_offset+15 && rot_y >= item_2_ingredient_2_y_offset && rot_y < item_2_ingredient_2_y_offset+15) begin
        case (item_2_id)
            2'b00: oled_data <= rice_boiled[14-(rot_y-item_2_ingredient_2_y_offset)] [14-(rot_x-item_2_ingredient_2_x_offset)];
            2'b01: oled_data <= cross[14-(rot_y-item_2_ingredient_2_y_offset)][14-(rot_x-item_2_ingredient_2_x_offset)];
            2'b10: oled_data <= cross[14-(rot_y-item_2_ingredient_2_y_offset)][14-(rot_x-item_2_ingredient_2_x_offset)];
            2'b11: oled_data <= rice_boiled[14-(rot_y-item_2_ingredient_2_y_offset)][14-(rot_x-item_2_ingredient_2_x_offset)];
        endcase
    end


    else if (rot_x >= item_3_ingredient_1_x_offset && rot_x < item_3_ingredient_1_x_offset+15 && rot_y >= item_3_ingredient_1_y_offset && rot_y < item_3_ingredient_1_y_offset+15) begin
        case (item_3_id)
            2'b00: oled_data <= chicken_boiled_chopped[14-(rot_y-item_3_ingredient_1_y_offset)][14-(rot_x-item_3_ingredient_1_x_offset)];
            2'b01: oled_data <= onion_boiled[14-(rot_y-item_3_ingredient_1_y_offset)][14-(rot_x-item_3_ingredient_1_x_offset)];
            2'b10: oled_data <= tomato_boiled[14-(rot_y-item_3_ingredient_1_y_offset)][14-(rot_x-item_3_ingredient_1_x_offset)];
            2'b11: oled_data <= tomato_boiled[14-(rot_y-item_3_ingredient_1_y_offset)][14-(rot_x-item_3_ingredient_1_x_offset)];
        endcase
    end

    else if (rot_x >= item_3_ingredient_2_x_offset && rot_x < item_3_ingredient_2_x_offset+15 && rot_y >= item_3_ingredient_2_y_offset && rot_y < item_3_ingredient_2_y_offset+15) begin
        case (item_3_id)
            2'b00: oled_data <= rice_boiled[14-(rot_y-item_3_ingredient_2_y_offset)][14-(rot_x-item_3_ingredient_2_x_offset)];
            2'b01: oled_data <= cross[14-(rot_y-item_3_ingredient_2_y_offset)][14-(rot_x-item_3_ingredient_2_x_offset)];
            2'b10: oled_data <= cross[14-(rot_y-item_3_ingredient_2_y_offset)][14-(rot_x-item_3_ingredient_2_x_offset)];
            2'b11: oled_data <= rice_boiled[14-(rot_y-item_3_ingredient_2_y_offset)][14-(rot_x-item_3_ingredient_2_x_offset)];
        endcase
    end

    else begin
        oled_data <= 0;
    end
end

endmodule


