module drawServe #(
    parameter [6:0] SERVE_TOP_LEFT_X = 0,
    parameter [6:0] SERVE_TOP_LEFT_Y = 0
)(
    input clk,
    input [6:0] x,
    input [6:0] y,
    output reg [15:0] oled_data
    );
    
    reg [15:0] serve1 [0:14][0:14];
    reg [15:0] serve2 [0:14][0:14];
    reg [15:0] serve3 [0:14][0:14];
    
    reg [6:0] x_idx;
    reg [6:0] y_idx;
    
    reg [1:0] state = 2'b00;
    
    wire slow_clock;
    reg prev_slow_clock = 0;
    wire frame_tick;
    
    flexible_clock frame_timer (
        .CLOCK(clk),
        .n(25_000_000),
        .SLOW_CLOCK(slow_clock)
    );
    
    // Rising edge detection
    assign frame_tick = (slow_clock == 1 && prev_slow_clock == 0);
    
    initial begin
    
        serve1[0][0] = 16'b11111_111110_11111;
    serve1[0][1] = 16'b11111_111110_11111;
    serve1[0][2] = 16'b11111_111110_11111;
    serve1[0][3] = 16'b11111_111110_11111;
    serve1[0][4] = 16'b11111_111110_11111;
    serve1[0][5] = 16'b11111_111110_11111;
    serve1[0][6] = 16'b11111_111110_11111;
    serve1[0][7] = 16'b11111_111110_11111;
    serve1[0][8] = 16'b11111_111110_11111;
    serve1[0][9] = 16'b11111_111110_11111;
    serve1[0][10] = 16'b11111_111110_11111;
    serve1[0][11] = 16'b11111_111110_11111;
    serve1[0][12] = 16'b11111_111110_11111;
    serve1[0][13] = 16'b11111_111110_11111;
    serve1[0][14] = 16'b11111_111110_11111;
    serve1[1][0] = 16'b11111_111110_11111;
    serve1[1][1] = 16'b00111_001111_00111;
    serve1[1][2] = 16'b00111_001111_00111;
    serve1[1][3] = 16'b00111_001111_00111;
    serve1[1][4] = 16'b00111_001111_00111;
    serve1[1][5] = 16'b00111_001111_00111;
    serve1[1][6] = 16'b00111_001111_00111;
    serve1[1][7] = 16'b00111_001111_00111;
    serve1[1][8] = 16'b00111_001111_00111;
    serve1[1][9] = 16'b00111_001111_00111;
    serve1[1][10] = 16'b00111_001111_00111;
    serve1[1][11] = 16'b00111_001111_00111;
    serve1[1][12] = 16'b00111_001111_00111;
    serve1[1][13] = 16'b00111_001111_00111;
    serve1[1][14] = 16'b11111_111110_11111;
    serve1[2][0] = 16'b11111_111110_11111;
    serve1[2][1] = 16'b00111_001111_00111;
    serve1[2][2] = 16'b00111_001111_00111;
    serve1[2][3] = 16'b00111_001111_00111;
    serve1[2][4] = 16'b00111_001111_00111;
    serve1[2][5] = 16'b00111_001111_00111;
    serve1[2][6] = 16'b00111_001111_00111;
    serve1[2][7] = 16'b00111_001111_00111;
    serve1[2][8] = 16'b00111_001111_00111;
    serve1[2][9] = 16'b00111_001111_00111;
    serve1[2][10] = 16'b00111_001111_00111;
    serve1[2][11] = 16'b00111_001111_00111;
    serve1[2][12] = 16'b00111_001111_00111;
    serve1[2][13] = 16'b00111_001111_00111;
    serve1[2][14] = 16'b11111_111110_11111;
    serve1[3][0] = 16'b11111_111110_11111;
    serve1[3][1] = 16'b00111_001111_00111;
    serve1[3][2] = 16'b01111_011111_01111;
    serve1[3][3] = 16'b01111_011111_01111;
    serve1[3][4] = 16'b01111_011111_01111;
    serve1[3][5] = 16'b01111_011111_01111;
    serve1[3][6] = 16'b01111_011111_01111;
    serve1[3][7] = 16'b01111_011111_01111;
    serve1[3][8] = 16'b01111_011111_01111;
    serve1[3][9] = 16'b01111_011111_01111;
    serve1[3][10] = 16'b01111_011111_01111;
    serve1[3][11] = 16'b01111_011111_01111;
    serve1[3][12] = 16'b01111_011111_01111;
    serve1[3][13] = 16'b00111_001111_00111;
    serve1[3][14] = 16'b11111_111110_11111;
    serve1[4][0] = 16'b11111_111110_11111;
    serve1[4][1] = 16'b00111_001111_00111;
    serve1[4][2] = 16'b00111_001111_00111;
    serve1[4][3] = 16'b01111_011111_01111;
    serve1[4][4] = 16'b01111_011111_01111;
    serve1[4][5] = 16'b01111_011111_01111;
    serve1[4][6] = 16'b01111_011111_01111;
    serve1[4][7] = 16'b01111_011111_01111;
    serve1[4][8] = 16'b01111_011111_01111;
    serve1[4][9] = 16'b01111_011111_01111;
    serve1[4][10] = 16'b01111_011111_01111;
    serve1[4][11] = 16'b01111_011111_01111;
    serve1[4][12] = 16'b00111_001111_00111;
    serve1[4][13] = 16'b00111_001111_00111;
    serve1[4][14] = 16'b11111_111110_11111;
    serve1[5][0] = 16'b11111_111110_11111;
    serve1[5][1] = 16'b00111_001111_00111;
    serve1[5][2] = 16'b00111_001111_00111;
    serve1[5][3] = 16'b00111_001111_00111;
    serve1[5][4] = 16'b01111_011111_01111;
    serve1[5][5] = 16'b01111_011111_01111;
    serve1[5][6] = 16'b01111_011111_01111;
    serve1[5][7] = 16'b01111_011111_01111;
    serve1[5][8] = 16'b01111_011111_01111;
    serve1[5][9] = 16'b01111_011111_01111;
    serve1[5][10] = 16'b01111_011111_01111;
    serve1[5][11] = 16'b00111_001111_00111;
    serve1[5][12] = 16'b00111_001111_00111;
    serve1[5][13] = 16'b00111_001111_00111;
    serve1[5][14] = 16'b11111_111110_11111;
    serve1[6][0] = 16'b11111_111110_11111;
    serve1[6][1] = 16'b00111_001111_00111;
    serve1[6][2] = 16'b00111_001111_00111;
    serve1[6][3] = 16'b00111_001111_00111;
    serve1[6][4] = 16'b00111_001111_00111;
    serve1[6][5] = 16'b01111_011111_01111;
    serve1[6][6] = 16'b01111_011111_01111;
    serve1[6][7] = 16'b01111_011111_01111;
    serve1[6][8] = 16'b01111_011111_01111;
    serve1[6][9] = 16'b01111_011111_01111;
    serve1[6][10] = 16'b00111_001111_00111;
    serve1[6][11] = 16'b00111_001111_00111;
    serve1[6][12] = 16'b00111_001111_00111;
    serve1[6][13] = 16'b00111_001111_00111;
    serve1[6][14] = 16'b11111_111110_11111;
    serve1[7][0] = 16'b11111_111110_11111;
    serve1[7][1] = 16'b00111_001111_00111;
    serve1[7][2] = 16'b00111_001111_00111;
    serve1[7][3] = 16'b00111_001111_00111;
    serve1[7][4] = 16'b00111_001111_00111;
    serve1[7][5] = 16'b00111_001111_00111;
    serve1[7][6] = 16'b01111_011111_01111;
    serve1[7][7] = 16'b01111_011111_01111;
    serve1[7][8] = 16'b01111_011111_01111;
    serve1[7][9] = 16'b00111_001111_00111;
    serve1[7][10] = 16'b00111_001111_00111;
    serve1[7][11] = 16'b00111_001111_00111;
    serve1[7][12] = 16'b00111_001111_00111;
    serve1[7][13] = 16'b00111_001111_00111;
    serve1[7][14] = 16'b11111_111110_11111;
    serve1[8][0] = 16'b11111_111110_11111;
    serve1[8][1] = 16'b00111_001111_00111;
    serve1[8][2] = 16'b00111_001111_00111;
    serve1[8][3] = 16'b00111_001111_00111;
    serve1[8][4] = 16'b00111_001111_00111;
    serve1[8][5] = 16'b00111_001111_00111;
    serve1[8][6] = 16'b00111_001111_00111;
    serve1[8][7] = 16'b01111_011111_01111;
    serve1[8][8] = 16'b00111_001111_00111;
    serve1[8][9] = 16'b00111_001111_00111;
    serve1[8][10] = 16'b00111_001111_00111;
    serve1[8][11] = 16'b00111_001111_00111;
    serve1[8][12] = 16'b00111_001111_00111;
    serve1[8][13] = 16'b00111_001111_00111;
    serve1[8][14] = 16'b11111_111110_11111;
    serve1[9][0] = 16'b11111_111110_11111;
    serve1[9][1] = 16'b00111_001111_00111;
    serve1[9][2] = 16'b00111_001111_00111;
    serve1[9][3] = 16'b00111_001111_00111;
    serve1[9][4] = 16'b00111_001111_00111;
    serve1[9][5] = 16'b00111_001111_00111;
    serve1[9][6] = 16'b00111_001111_00111;
    serve1[9][7] = 16'b00111_001111_00111;
    serve1[9][8] = 16'b00111_001111_00111;
    serve1[9][9] = 16'b00111_001111_00111;
    serve1[9][10] = 16'b00111_001111_00111;
    serve1[9][11] = 16'b00111_001111_00111;
    serve1[9][12] = 16'b00111_001111_00111;
    serve1[9][13] = 16'b00111_001111_00111;
    serve1[9][14] = 16'b11111_111110_11111;
    serve1[10][0] = 16'b11111_111110_11111;
    serve1[10][1] = 16'b00111_001111_00111;
    serve1[10][2] = 16'b00111_001111_00111;
    serve1[10][3] = 16'b00111_001111_00111;
    serve1[10][4] = 16'b00111_001111_00111;
    serve1[10][5] = 16'b00111_001111_00111;
    serve1[10][6] = 16'b00111_001111_00111;
    serve1[10][7] = 16'b00111_001111_00111;
    serve1[10][8] = 16'b00111_001111_00111;
    serve1[10][9] = 16'b00111_001111_00111;
    serve1[10][10] = 16'b00111_001111_00111;
    serve1[10][11] = 16'b00111_001111_00111;
    serve1[10][12] = 16'b00111_001111_00111;
    serve1[10][13] = 16'b00111_001111_00111;
    serve1[10][14] = 16'b11111_111110_11111;
    serve1[11][0] = 16'b11111_111110_11111;
    serve1[11][1] = 16'b00111_001111_00111;
    serve1[11][2] = 16'b00111_001111_00111;
    serve1[11][3] = 16'b00111_001111_00111;
    serve1[11][4] = 16'b00111_001111_00111;
    serve1[11][5] = 16'b00111_001111_00111;
    serve1[11][6] = 16'b00111_001111_00111;
    serve1[11][7] = 16'b00111_001111_00111;
    serve1[11][8] = 16'b00111_001111_00111;
    serve1[11][9] = 16'b00111_001111_00111;
    serve1[11][10] = 16'b00111_001111_00111;
    serve1[11][11] = 16'b00111_001111_00111;
    serve1[11][12] = 16'b00111_001111_00111;
    serve1[11][13] = 16'b00111_001111_00111;
    serve1[11][14] = 16'b11111_111110_11111;
    serve1[12][0] = 16'b11111_111110_11111;
    serve1[12][1] = 16'b00111_001111_00111;
    serve1[12][2] = 16'b00111_001111_00111;
    serve1[12][3] = 16'b00111_001111_00111;
    serve1[12][4] = 16'b00111_001111_00111;
    serve1[12][5] = 16'b00111_001111_00111;
    serve1[12][6] = 16'b00111_001111_00111;
    serve1[12][7] = 16'b00111_001111_00111;
    serve1[12][8] = 16'b00111_001111_00111;
    serve1[12][9] = 16'b00111_001111_00111;
    serve1[12][10] = 16'b00111_001111_00111;
    serve1[12][11] = 16'b00111_001111_00111;
    serve1[12][12] = 16'b00111_001111_00111;
    serve1[12][13] = 16'b00111_001111_00111;
    serve1[12][14] = 16'b11111_111110_11111;
    serve1[13][0] = 16'b11111_111110_11111;
    serve1[13][1] = 16'b00111_001111_00111;
    serve1[13][2] = 16'b00111_001111_00111;
    serve1[13][3] = 16'b00111_001111_00111;
    serve1[13][4] = 16'b00111_001111_00111;
    serve1[13][5] = 16'b00111_001111_00111;
    serve1[13][6] = 16'b00111_001111_00111;
    serve1[13][7] = 16'b00111_001111_00111;
    serve1[13][8] = 16'b00111_001111_00111;
    serve1[13][9] = 16'b00111_001111_00111;
    serve1[13][10] = 16'b00111_001111_00111;
    serve1[13][11] = 16'b00111_001111_00111;
    serve1[13][12] = 16'b00111_001111_00111;
    serve1[13][13] = 16'b00111_001111_00111;
    serve1[13][14] = 16'b11111_111110_11111;
    serve1[14][0] = 16'b11111_111110_11111;
    serve1[14][1] = 16'b11111_111110_11111;
    serve1[14][2] = 16'b11111_111110_11111;
    serve1[14][3] = 16'b11111_111110_11111;
    serve1[14][4] = 16'b11111_111110_11111;
    serve1[14][5] = 16'b11111_111110_11111;
    serve1[14][6] = 16'b11111_111110_11111;
    serve1[14][7] = 16'b11111_111110_11111;
    serve1[14][8] = 16'b11111_111110_11111;
    serve1[14][9] = 16'b11111_111110_11111;
    serve1[14][10] = 16'b11111_111110_11111;
    serve1[14][11] = 16'b11111_111110_11111;
    serve1[14][12] = 16'b11111_111110_11111;
    serve1[14][13] = 16'b11111_111110_11111;
    serve1[14][14] = 16'b11111_111110_11111;

    serve2[0][0] = 16'b11111_111110_11111;
    serve2[0][1] = 16'b11111_111110_11111;
    serve2[0][2] = 16'b11111_111110_11111;
    serve2[0][3] = 16'b11111_111110_11111;
    serve2[0][4] = 16'b11111_111110_11111;
    serve2[0][5] = 16'b11111_111110_11111;
    serve2[0][6] = 16'b11111_111110_11111;
    serve2[0][7] = 16'b11111_111110_11111;
    serve2[0][8] = 16'b11111_111110_11111;
    serve2[0][9] = 16'b11111_111110_11111;
    serve2[0][10] = 16'b11111_111110_11111;
    serve2[0][11] = 16'b11111_111110_11111;
    serve2[0][12] = 16'b11111_111110_11111;
    serve2[0][13] = 16'b11111_111110_11111;
    serve2[0][14] = 16'b11111_111110_11111;
    serve2[1][0] = 16'b11111_111110_11111;
    serve2[1][1] = 16'b00111_001111_00111;
    serve2[1][2] = 16'b00111_001111_00111;
    serve2[1][3] = 16'b00111_001111_00111;
    serve2[1][4] = 16'b00111_001111_00111;
    serve2[1][5] = 16'b00111_001111_00111;
    serve2[1][6] = 16'b00111_001111_00111;
    serve2[1][7] = 16'b00111_001111_00111;
    serve2[1][8] = 16'b00111_001111_00111;
    serve2[1][9] = 16'b00111_001111_00111;
    serve2[1][10] = 16'b00111_001111_00111;
    serve2[1][11] = 16'b00111_001111_00111;
    serve2[1][12] = 16'b00111_001111_00111;
    serve2[1][13] = 16'b00111_001111_00111;
    serve2[1][14] = 16'b11111_111110_11111;
    serve2[2][0] = 16'b11111_111110_11111;
    serve2[2][1] = 16'b00111_001111_00111;
    serve2[2][2] = 16'b00111_001111_00111;
    serve2[2][3] = 16'b00111_001111_00111;
    serve2[2][4] = 16'b00111_001111_00111;
    serve2[2][5] = 16'b00111_001111_00111;
    serve2[2][6] = 16'b00111_001111_00111;
    serve2[2][7] = 16'b00111_001111_00111;
    serve2[2][8] = 16'b00111_001111_00111;
    serve2[2][9] = 16'b00111_001111_00111;
    serve2[2][10] = 16'b00111_001111_00111;
    serve2[2][11] = 16'b00111_001111_00111;
    serve2[2][12] = 16'b00111_001111_00111;
    serve2[2][13] = 16'b00111_001111_00111;
    serve2[2][14] = 16'b11111_111110_11111;
    serve2[3][0] = 16'b11111_111110_11111;
    serve2[3][1] = 16'b00111_001111_00111;
    serve2[3][2] = 16'b00111_001111_00111;
    serve2[3][3] = 16'b00111_001111_00111;
    serve2[3][4] = 16'b00111_001111_00111;
    serve2[3][5] = 16'b00111_001111_00111;
    serve2[3][6] = 16'b00111_001111_00111;
    serve2[3][7] = 16'b00111_001111_00111;
    serve2[3][8] = 16'b00111_001111_00111;
    serve2[3][9] = 16'b00111_001111_00111;
    serve2[3][10] = 16'b00111_001111_00111;
    serve2[3][11] = 16'b00111_001111_00111;
    serve2[3][12] = 16'b00111_001111_00111;
    serve2[3][13] = 16'b00111_001111_00111;
    serve2[3][14] = 16'b11111_111110_11111;
    serve2[4][0] = 16'b11111_111110_11111;
    serve2[4][1] = 16'b00111_001111_00111;
    serve2[4][2] = 16'b00111_001111_00111;
    serve2[4][3] = 16'b00111_001111_00111;
    serve2[4][4] = 16'b00111_001111_00111;
    serve2[4][5] = 16'b00111_001111_00111;
    serve2[4][6] = 16'b00111_001111_00111;
    serve2[4][7] = 16'b00111_001111_00111;
    serve2[4][8] = 16'b00111_001111_00111;
    serve2[4][9] = 16'b00111_001111_00111;
    serve2[4][10] = 16'b00111_001111_00111;
    serve2[4][11] = 16'b00111_001111_00111;
    serve2[4][12] = 16'b00111_001111_00111;
    serve2[4][13] = 16'b00111_001111_00111;
    serve2[4][14] = 16'b11111_111110_11111;
    serve2[5][0] = 16'b11111_111110_11111;
    serve2[5][1] = 16'b00111_001111_00111;
    serve2[5][2] = 16'b01111_011111_01111;
    serve2[5][3] = 16'b01111_011111_01111;
    serve2[5][4] = 16'b01111_011111_01111;
    serve2[5][5] = 16'b01111_011111_01111;
    serve2[5][6] = 16'b01111_011111_01111;
    serve2[5][7] = 16'b01111_011111_01111;
    serve2[5][8] = 16'b01111_011111_01111;
    serve2[5][9] = 16'b01111_011111_01111;
    serve2[5][10] = 16'b01111_011111_01111;
    serve2[5][11] = 16'b01111_011111_01111;
    serve2[5][12] = 16'b01111_011111_01111;
    serve2[5][13] = 16'b00111_001111_00111;
    serve2[5][14] = 16'b11111_111110_11111;
    serve2[6][0] = 16'b11111_111110_11111;
    serve2[6][1] = 16'b00111_001111_00111;
    serve2[6][2] = 16'b00111_001111_00111;
    serve2[6][3] = 16'b01111_011111_01111;
    serve2[6][4] = 16'b01111_011111_01111;
    serve2[6][5] = 16'b01111_011111_01111;
    serve2[6][6] = 16'b01111_011111_01111;
    serve2[6][7] = 16'b01111_011111_01111;
    serve2[6][8] = 16'b01111_011111_01111;
    serve2[6][9] = 16'b01111_011111_01111;
    serve2[6][10] = 16'b01111_011111_01111;
    serve2[6][11] = 16'b01111_011111_01111;
    serve2[6][12] = 16'b00111_001111_00111;
    serve2[6][13] = 16'b00111_001111_00111;
    serve2[6][14] = 16'b11111_111110_11111;
    serve2[7][0] = 16'b11111_111110_11111;
    serve2[7][1] = 16'b00111_001111_00111;
    serve2[7][2] = 16'b00111_001111_00111;
    serve2[7][3] = 16'b00111_001111_00111;
    serve2[7][4] = 16'b01111_011111_01111;
    serve2[7][5] = 16'b01111_011111_01111;
    serve2[7][6] = 16'b01111_011111_01111;
    serve2[7][7] = 16'b01111_011111_01111;
    serve2[7][8] = 16'b01111_011111_01111;
    serve2[7][9] = 16'b01111_011111_01111;
    serve2[7][10] = 16'b01111_011111_01111;
    serve2[7][11] = 16'b00111_001111_00111;
    serve2[7][12] = 16'b00111_001111_00111;
    serve2[7][13] = 16'b00111_001111_00111;
    serve2[7][14] = 16'b11111_111110_11111;
    serve2[8][0] = 16'b11111_111110_11111;
    serve2[8][1] = 16'b00111_001111_00111;
    serve2[8][2] = 16'b00111_001111_00111;
    serve2[8][3] = 16'b00111_001111_00111;
    serve2[8][4] = 16'b00111_001111_00111;
    serve2[8][5] = 16'b01111_011111_01111;
    serve2[8][6] = 16'b01111_011111_01111;
    serve2[8][7] = 16'b01111_011111_01111;
    serve2[8][8] = 16'b01111_011111_01111;
    serve2[8][9] = 16'b01111_011111_01111;
    serve2[8][10] = 16'b00111_001111_00111;
    serve2[8][11] = 16'b00111_001111_00111;
    serve2[8][12] = 16'b00111_001111_00111;
    serve2[8][13] = 16'b00111_001111_00111;
    serve2[8][14] = 16'b11111_111110_11111;
    serve2[9][0] = 16'b11111_111110_11111;
    serve2[9][1] = 16'b00111_001111_00111;
    serve2[9][2] = 16'b00111_001111_00111;
    serve2[9][3] = 16'b00111_001111_00111;
    serve2[9][4] = 16'b00111_001111_00111;
    serve2[9][5] = 16'b00111_001111_00111;
    serve2[9][6] = 16'b01111_011111_01111;
    serve2[9][7] = 16'b01111_011111_01111;
    serve2[9][8] = 16'b01111_011111_01111;
    serve2[9][9] = 16'b00111_001111_00111;
    serve2[9][10] = 16'b00111_001111_00111;
    serve2[9][11] = 16'b00111_001111_00111;
    serve2[9][12] = 16'b00111_001111_00111;
    serve2[9][13] = 16'b00111_001111_00111;
    serve2[9][14] = 16'b11111_111110_11111;
    serve2[10][0] = 16'b11111_111110_11111;
    serve2[10][1] = 16'b00111_001111_00111;
    serve2[10][2] = 16'b00111_001111_00111;
    serve2[10][3] = 16'b00111_001111_00111;
    serve2[10][4] = 16'b00111_001111_00111;
    serve2[10][5] = 16'b00111_001111_00111;
    serve2[10][6] = 16'b00111_001111_00111;
    serve2[10][7] = 16'b01111_011111_01111;
    serve2[10][8] = 16'b00111_001111_00111;
    serve2[10][9] = 16'b00111_001111_00111;
    serve2[10][10] = 16'b00111_001111_00111;
    serve2[10][11] = 16'b00111_001111_00111;
    serve2[10][12] = 16'b00111_001111_00111;
    serve2[10][13] = 16'b00111_001111_00111;
    serve2[10][14] = 16'b11111_111110_11111;
    serve2[11][0] = 16'b11111_111110_11111;
    serve2[11][1] = 16'b00111_001111_00111;
    serve2[11][2] = 16'b00111_001111_00111;
    serve2[11][3] = 16'b00111_001111_00111;
    serve2[11][4] = 16'b00111_001111_00111;
    serve2[11][5] = 16'b00111_001111_00111;
    serve2[11][6] = 16'b00111_001111_00111;
    serve2[11][7] = 16'b00111_001111_00111;
    serve2[11][8] = 16'b00111_001111_00111;
    serve2[11][9] = 16'b00111_001111_00111;
    serve2[11][10] = 16'b00111_001111_00111;
    serve2[11][11] = 16'b00111_001111_00111;
    serve2[11][12] = 16'b00111_001111_00111;
    serve2[11][13] = 16'b00111_001111_00111;
    serve2[11][14] = 16'b11111_111110_11111;
    serve2[12][0] = 16'b11111_111110_11111;
    serve2[12][1] = 16'b00111_001111_00111;
    serve2[12][2] = 16'b00111_001111_00111;
    serve2[12][3] = 16'b00111_001111_00111;
    serve2[12][4] = 16'b00111_001111_00111;
    serve2[12][5] = 16'b00111_001111_00111;
    serve2[12][6] = 16'b00111_001111_00111;
    serve2[12][7] = 16'b00111_001111_00111;
    serve2[12][8] = 16'b00111_001111_00111;
    serve2[12][9] = 16'b00111_001111_00111;
    serve2[12][10] = 16'b00111_001111_00111;
    serve2[12][11] = 16'b00111_001111_00111;
    serve2[12][12] = 16'b00111_001111_00111;
    serve2[12][13] = 16'b00111_001111_00111;
    serve2[12][14] = 16'b11111_111110_11111;
    serve2[13][0] = 16'b11111_111110_11111;
    serve2[13][1] = 16'b00111_001111_00111;
    serve2[13][2] = 16'b00111_001111_00111;
    serve2[13][3] = 16'b00111_001111_00111;
    serve2[13][4] = 16'b00111_001111_00111;
    serve2[13][5] = 16'b00111_001111_00111;
    serve2[13][6] = 16'b00111_001111_00111;
    serve2[13][7] = 16'b00111_001111_00111;
    serve2[13][8] = 16'b00111_001111_00111;
    serve2[13][9] = 16'b00111_001111_00111;
    serve2[13][10] = 16'b00111_001111_00111;
    serve2[13][11] = 16'b00111_001111_00111;
    serve2[13][12] = 16'b00111_001111_00111;
    serve2[13][13] = 16'b00111_001111_00111;
    serve2[13][14] = 16'b11111_111110_11111;
    serve2[14][0] = 16'b11111_111110_11111;
    serve2[14][1] = 16'b11111_111110_11111;
    serve2[14][2] = 16'b11111_111110_11111;
    serve2[14][3] = 16'b11111_111110_11111;
    serve2[14][4] = 16'b11111_111110_11111;
    serve2[14][5] = 16'b11111_111110_11111;
    serve2[14][6] = 16'b11111_111110_11111;
    serve2[14][7] = 16'b11111_111110_11111;
    serve2[14][8] = 16'b11111_111110_11111;
    serve2[14][9] = 16'b11111_111110_11111;
    serve2[14][10] = 16'b11111_111110_11111;
    serve2[14][11] = 16'b11111_111110_11111;
    serve2[14][12] = 16'b11111_111110_11111;
    serve2[14][13] = 16'b11111_111110_11111;
    serve2[14][14] = 16'b11111_111110_11111;
    
    serve3[0][0] = 16'b11111_111110_11111;
    serve3[0][1] = 16'b11111_111110_11111;
    serve3[0][2] = 16'b11111_111110_11111;
    serve3[0][3] = 16'b11111_111110_11111;
    serve3[0][4] = 16'b11111_111110_11111;
    serve3[0][5] = 16'b11111_111110_11111;
    serve3[0][6] = 16'b11111_111110_11111;
    serve3[0][7] = 16'b11111_111110_11111;
    serve3[0][8] = 16'b11111_111110_11111;
    serve3[0][9] = 16'b11111_111110_11111;
    serve3[0][10] = 16'b11111_111110_11111;
    serve3[0][11] = 16'b11111_111110_11111;
    serve3[0][12] = 16'b11111_111110_11111;
    serve3[0][13] = 16'b11111_111110_11111;
    serve3[0][14] = 16'b11111_111110_11111;
    serve3[1][0] = 16'b11111_111110_11111;
    serve3[1][1] = 16'b00111_001111_00111;
    serve3[1][2] = 16'b00111_001111_00111;
    serve3[1][3] = 16'b00111_001111_00111;
    serve3[1][4] = 16'b00111_001111_00111;
    serve3[1][5] = 16'b00111_001111_00111;
    serve3[1][6] = 16'b00111_001111_00111;
    serve3[1][7] = 16'b00111_001111_00111;
    serve3[1][8] = 16'b00111_001111_00111;
    serve3[1][9] = 16'b00111_001111_00111;
    serve3[1][10] = 16'b00111_001111_00111;
    serve3[1][11] = 16'b00111_001111_00111;
    serve3[1][12] = 16'b00111_001111_00111;
    serve3[1][13] = 16'b00111_001111_00111;
    serve3[1][14] = 16'b11111_111110_11111;
    serve3[2][0] = 16'b11111_111110_11111;
    serve3[2][1] = 16'b00111_001111_00111;
    serve3[2][2] = 16'b00111_001111_00111;
    serve3[2][3] = 16'b00111_001111_00111;
    serve3[2][4] = 16'b00111_001111_00111;
    serve3[2][5] = 16'b00111_001111_00111;
    serve3[2][6] = 16'b00111_001111_00111;
    serve3[2][7] = 16'b00111_001111_00111;
    serve3[2][8] = 16'b00111_001111_00111;
    serve3[2][9] = 16'b00111_001111_00111;
    serve3[2][10] = 16'b00111_001111_00111;
    serve3[2][11] = 16'b00111_001111_00111;
    serve3[2][12] = 16'b00111_001111_00111;
    serve3[2][13] = 16'b00111_001111_00111;
    serve3[2][14] = 16'b11111_111110_11111;
    serve3[3][0] = 16'b11111_111110_11111;
    serve3[3][1] = 16'b00111_001111_00111;
    serve3[3][2] = 16'b00111_001111_00111;
    serve3[3][3] = 16'b00111_001111_00111;
    serve3[3][4] = 16'b00111_001111_00111;
    serve3[3][5] = 16'b00111_001111_00111;
    serve3[3][6] = 16'b00111_001111_00111;
    serve3[3][7] = 16'b00111_001111_00111;
    serve3[3][8] = 16'b00111_001111_00111;
    serve3[3][9] = 16'b00111_001111_00111;
    serve3[3][10] = 16'b00111_001111_00111;
    serve3[3][11] = 16'b00111_001111_00111;
    serve3[3][12] = 16'b00111_001111_00111;
    serve3[3][13] = 16'b00111_001111_00111;
    serve3[3][14] = 16'b11111_111110_11111;
    serve3[4][0] = 16'b11111_111110_11111;
    serve3[4][1] = 16'b00111_001111_00111;
    serve3[4][2] = 16'b00111_001111_00111;
    serve3[4][3] = 16'b00111_001111_00111;
    serve3[4][4] = 16'b00111_001111_00111;
    serve3[4][5] = 16'b00111_001111_00111;
    serve3[4][6] = 16'b00111_001111_00111;
    serve3[4][7] = 16'b00111_001111_00111;
    serve3[4][8] = 16'b00111_001111_00111;
    serve3[4][9] = 16'b00111_001111_00111;
    serve3[4][10] = 16'b00111_001111_00111;
    serve3[4][11] = 16'b00111_001111_00111;
    serve3[4][12] = 16'b00111_001111_00111;
    serve3[4][13] = 16'b00111_001111_00111;
    serve3[4][14] = 16'b11111_111110_11111;
    serve3[5][0] = 16'b11111_111110_11111;
    serve3[5][1] = 16'b00111_001111_00111;
    serve3[5][2] = 16'b00111_001111_00111;
    serve3[5][3] = 16'b00111_001111_00111;
    serve3[5][4] = 16'b00111_001111_00111;
    serve3[5][5] = 16'b00111_001111_00111;
    serve3[5][6] = 16'b00111_001111_00111;
    serve3[5][7] = 16'b00111_001111_00111;
    serve3[5][8] = 16'b00111_001111_00111;
    serve3[5][9] = 16'b00111_001111_00111;
    serve3[5][10] = 16'b00111_001111_00111;
    serve3[5][11] = 16'b00111_001111_00111;
    serve3[5][12] = 16'b00111_001111_00111;
    serve3[5][13] = 16'b00111_001111_00111;
    serve3[5][14] = 16'b11111_111110_11111;
    serve3[6][0] = 16'b11111_111110_11111;
    serve3[6][1] = 16'b00111_001111_00111;
    serve3[6][2] = 16'b00111_001111_00111;
    serve3[6][3] = 16'b00111_001111_00111;
    serve3[6][4] = 16'b00111_001111_00111;
    serve3[6][5] = 16'b00111_001111_00111;
    serve3[6][6] = 16'b00111_001111_00111;
    serve3[6][7] = 16'b00111_001111_00111;
    serve3[6][8] = 16'b00111_001111_00111;
    serve3[6][9] = 16'b00111_001111_00111;
    serve3[6][10] = 16'b00111_001111_00111;
    serve3[6][11] = 16'b00111_001111_00111;
    serve3[6][12] = 16'b00111_001111_00111;
    serve3[6][13] = 16'b00111_001111_00111;
    serve3[6][14] = 16'b11111_111110_11111;
    serve3[7][0] = 16'b11111_111110_11111;
    serve3[7][1] = 16'b00111_001111_00111;
    serve3[7][2] = 16'b01111_011111_01111;
    serve3[7][3] = 16'b01111_011111_01111;
    serve3[7][4] = 16'b01111_011111_01111;
    serve3[7][5] = 16'b01111_011111_01111;
    serve3[7][6] = 16'b01111_011111_01111;
    serve3[7][7] = 16'b01111_011111_01111;
    serve3[7][8] = 16'b01111_011111_01111;
    serve3[7][9] = 16'b01111_011111_01111;
    serve3[7][10] = 16'b01111_011111_01111;
    serve3[7][11] = 16'b01111_011111_01111;
    serve3[7][12] = 16'b01111_011111_01111;
    serve3[7][13] = 16'b00111_001111_00111;
    serve3[7][14] = 16'b11111_111110_11111;
    serve3[8][0] = 16'b11111_111110_11111;
    serve3[8][1] = 16'b00111_001111_00111;
    serve3[8][2] = 16'b00111_001111_00111;
    serve3[8][3] = 16'b01111_011111_01111;
    serve3[8][4] = 16'b01111_011111_01111;
    serve3[8][5] = 16'b01111_011111_01111;
    serve3[8][6] = 16'b01111_011111_01111;
    serve3[8][7] = 16'b01111_011111_01111;
    serve3[8][8] = 16'b01111_011111_01111;
    serve3[8][9] = 16'b01111_011111_01111;
    serve3[8][10] = 16'b01111_011111_01111;
    serve3[8][11] = 16'b01111_011111_01111;
    serve3[8][12] = 16'b00111_001111_00111;
    serve3[8][13] = 16'b00111_001111_00111;
    serve3[8][14] = 16'b11111_111110_11111;
    serve3[9][0] = 16'b11111_111110_11111;
    serve3[9][1] = 16'b00111_001111_00111;
    serve3[9][2] = 16'b00111_001111_00111;
    serve3[9][3] = 16'b00111_001111_00111;
    serve3[9][4] = 16'b01111_011111_01111;
    serve3[9][5] = 16'b01111_011111_01111;
    serve3[9][6] = 16'b01111_011111_01111;
    serve3[9][7] = 16'b01111_011111_01111;
    serve3[9][8] = 16'b01111_011111_01111;
    serve3[9][9] = 16'b01111_011111_01111;
    serve3[9][10] = 16'b01111_011111_01111;
    serve3[9][11] = 16'b00111_001111_00111;
    serve3[9][12] = 16'b00111_001111_00111;
    serve3[9][13] = 16'b00111_001111_00111;
    serve3[9][14] = 16'b11111_111110_11111;
    serve3[10][0] = 16'b11111_111110_11111;
    serve3[10][1] = 16'b00111_001111_00111;
    serve3[10][2] = 16'b00111_001111_00111;
    serve3[10][3] = 16'b00111_001111_00111;
    serve3[10][4] = 16'b00111_001111_00111;
    serve3[10][5] = 16'b01111_011111_01111;
    serve3[10][6] = 16'b01111_011111_01111;
    serve3[10][7] = 16'b01111_011111_01111;
    serve3[10][8] = 16'b01111_011111_01111;
    serve3[10][9] = 16'b01111_011111_01111;
    serve3[10][10] = 16'b00111_001111_00111;
    serve3[10][11] = 16'b00111_001111_00111;
    serve3[10][12] = 16'b00111_001111_00111;
    serve3[10][13] = 16'b00111_001111_00111;
    serve3[10][14] = 16'b11111_111110_11111;
    serve3[11][0] = 16'b11111_111110_11111;
    serve3[11][1] = 16'b00111_001111_00111;
    serve3[11][2] = 16'b00111_001111_00111;
    serve3[11][3] = 16'b00111_001111_00111;
    serve3[11][4] = 16'b00111_001111_00111;
    serve3[11][5] = 16'b00111_001111_00111;
    serve3[11][6] = 16'b01111_011111_01111;
    serve3[11][7] = 16'b01111_011111_01111;
    serve3[11][8] = 16'b01111_011111_01111;
    serve3[11][9] = 16'b00111_001111_00111;
    serve3[11][10] = 16'b00111_001111_00111;
    serve3[11][11] = 16'b00111_001111_00111;
    serve3[11][12] = 16'b00111_001111_00111;
    serve3[11][13] = 16'b00111_001111_00111;
    serve3[11][14] = 16'b11111_111110_11111;
    serve3[12][0] = 16'b11111_111110_11111;
    serve3[12][1] = 16'b00111_001111_00111;
    serve3[12][2] = 16'b00111_001111_00111;
    serve3[12][3] = 16'b00111_001111_00111;
    serve3[12][4] = 16'b00111_001111_00111;
    serve3[12][5] = 16'b00111_001111_00111;
    serve3[12][6] = 16'b00111_001111_00111;
    serve3[12][7] = 16'b01111_011111_01111;
    serve3[12][8] = 16'b00111_001111_00111;
    serve3[12][9] = 16'b00111_001111_00111;
    serve3[12][10] = 16'b00111_001111_00111;
    serve3[12][11] = 16'b00111_001111_00111;
    serve3[12][12] = 16'b00111_001111_00111;
    serve3[12][13] = 16'b00111_001111_00111;
    serve3[12][14] = 16'b11111_111110_11111;
    serve3[13][0] = 16'b11111_111110_11111;
    serve3[13][1] = 16'b00111_001111_00111;
    serve3[13][2] = 16'b00111_001111_00111;
    serve3[13][3] = 16'b00111_001111_00111;
    serve3[13][4] = 16'b00111_001111_00111;
    serve3[13][5] = 16'b00111_001111_00111;
    serve3[13][6] = 16'b00111_001111_00111;
    serve3[13][7] = 16'b00111_001111_00111;
    serve3[13][8] = 16'b00111_001111_00111;
    serve3[13][9] = 16'b00111_001111_00111;
    serve3[13][10] = 16'b00111_001111_00111;
    serve3[13][11] = 16'b00111_001111_00111;
    serve3[13][12] = 16'b00111_001111_00111;
    serve3[13][13] = 16'b00111_001111_00111;
    serve3[13][14] = 16'b11111_111110_11111;
    serve3[14][0] = 16'b11111_111110_11111;
    serve3[14][1] = 16'b11111_111110_11111;
    serve3[14][2] = 16'b11111_111110_11111;
    serve3[14][3] = 16'b11111_111110_11111;
    serve3[14][4] = 16'b11111_111110_11111;
    serve3[14][5] = 16'b11111_111110_11111;
    serve3[14][6] = 16'b11111_111110_11111;
    serve3[14][7] = 16'b11111_111110_11111;
    serve3[14][8] = 16'b11111_111110_11111;
    serve3[14][9] = 16'b11111_111110_11111;
    serve3[14][10] = 16'b11111_111110_11111;
    serve3[14][11] = 16'b11111_111110_11111;
    serve3[14][12] = 16'b11111_111110_11111;
    serve3[14][13] = 16'b11111_111110_11111;
    serve3[14][14] = 16'b11111_111110_11111;

    end
    
    always @(posedge clk) begin
        prev_slow_clock <= slow_clock;
        
        case (state)
            2'd0: if (frame_tick) state <= 2'd1;
            2'd1: if (frame_tick) state <= 2'd2;
            2'd2: if (frame_tick) state <= 2'd3;
            2'd3: if (frame_tick) state <= 2'd0;
        endcase
        
    end
    
    always @(*) begin
        x_idx = x - SERVE_TOP_LEFT_X;
        y_idx = y - SERVE_TOP_LEFT_Y;
        
        if (x_idx >= 0 && x_idx < 15 && y_idx >= 0 && y_idx < 15) begin
            case (state)
                2'd0: oled_data = serve1[y_idx][x_idx];
                2'd1: oled_data = serve2[y_idx][x_idx];
                2'd2: oled_data = serve3[y_idx][x_idx];
                2'd3: oled_data = serve2[y_idx][x_idx];
                default: oled_data = serve2[y_idx][x_idx];
            endcase
        end else begin
            oled_data = 0;
        end
        
    end
    
    
endmodule
