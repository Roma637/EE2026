`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08.04.2025 21:20:34
// Design Name: 
// Module Name: draw_chopper
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module draw_chopper #(
    parameter [6:0] CHOPPER_TOP_LEFT_X = 0,
    parameter [6:0] CHOPPER_TOP_LEFT_Y = 0
)(
    input clk,
    input chop_ready,
    input reset,
    input [7:0] x,
    input [6:0] y,
    output reg [15:0] oled_data
    );
    
    reg [15:0] chop_empty [0:14][0:14];
    reg [15:0] chop_full [0:14][0:14];
    
    reg [15:0] timing1 [0:14][0:14];
    reg [15:0] timing2 [0:14][0:14];
    reg [15:0] timing3 [0:14][0:14];
    reg [15:0] timing4 [0:14][0:14];
    reg [15:0] timing5 [0:14][0:14];
    reg [15:0] timing6 [0:14][0:14];
    reg [15:0] timing7 [0:14][0:14];
    reg [15:0] timing8 [0:14][0:14];
    reg [15:0] timing9 [0:14][0:14];
    
    reg [7:0] x_idx;
    reg [6:0] y_idx;
    
    // 00 - empty
    // 01 - clocks
    // 10 - full
    reg [3:0] state = 0;
    localparam IDLE = 0;
    localparam ANIM1 = 1;
    localparam ANIM2 = 2;
    localparam ANIM3 = 3;
    localparam ANIM4 = 4;
    localparam ANIM5 = 5;
    localparam ANIM6 = 6;
    localparam ANIM7 = 7;
    localparam ANIM8 = 8;
    localparam ANIM9 = 9;
    localparam FULL = 10;
    
    wire slow_clock;
    reg prev_slow_clock = 0;
    wire frame_tick;
    
    flexible_clock frame_timer (
        clk,
        25_000_000,
        slow_clock
    );
    
    // Rising edge detection
    assign frame_tick = (slow_clock == 1 && prev_slow_clock == 0);

    
//    flexible_clock #(25_000_000) frame_timer (
//        .clk(clk),
//        .enable(enable_clock),
//        .tick(frame_tick)
//    );
    
//    flexible_clock frame_timer(
//        .clk(clk),
//        .signal(frame_tick),
//        .n(12_500_000)
//    );
    
    initial begin
    
    state = 2'b0;

    timing1[0][0] = 16'b11111_111110_11111;
    timing1[0][1] = 16'b11111_111110_11111;
    timing1[0][2] = 16'b11111_111110_11111;
    timing1[0][3] = 16'b11111_111110_11111;
    timing1[0][4] = 16'b11111_111110_11111;
    timing1[0][5] = 16'b11111_111110_11111;
    timing1[0][6] = 16'b11111_111110_11111;
    timing1[0][7] = 16'b11111_111110_11111;
    timing1[0][8] = 16'b11111_111110_11111;
    timing1[0][9] = 16'b11111_111110_11111;
    timing1[0][10] = 16'b11111_111110_11111;
    timing1[0][11] = 16'b11111_111110_11111;
    timing1[0][12] = 16'b11111_111110_11111;
    timing1[0][13] = 16'b11111_111110_11111;
    timing1[0][14] = 16'b11111_111110_11111;
    timing1[1][0] = 16'b11111_111110_11111;
    timing1[1][1] = 16'b00000_000000_00000;
    timing1[1][2] = 16'b00000_000000_00000;
    timing1[1][3] = 16'b00000_000000_00000;
    timing1[1][4] = 16'b00000_000000_00000;
    timing1[1][5] = 16'b11111_101110_00000;
    timing1[1][6] = 16'b11111_101110_00000;
    timing1[1][7] = 16'b11111_101110_00000;
    timing1[1][8] = 16'b11111_101110_00000;
    timing1[1][9] = 16'b11111_101110_00000;
    timing1[1][10] = 16'b00000_000000_00000;
    timing1[1][11] = 16'b00000_000000_00000;
    timing1[1][12] = 16'b00000_000000_00000;
    timing1[1][13] = 16'b00000_000000_00000;
    timing1[1][14] = 16'b11111_111110_11111;
    timing1[2][0] = 16'b11111_111110_11111;
    timing1[2][1] = 16'b00000_000000_00000;
    timing1[2][2] = 16'b00000_000000_00000;
    timing1[2][3] = 16'b11111_101110_00000;
    timing1[2][4] = 16'b11111_101110_00000;
    timing1[2][5] = 16'b11001_100100_00000;
    timing1[2][6] = 16'b11001_100100_00000;
    timing1[2][7] = 16'b11001_100100_00000;
    timing1[2][8] = 16'b11001_100100_00000;
    timing1[2][9] = 16'b11001_100100_00000;
    timing1[2][10] = 16'b11111_101110_00000;
    timing1[2][11] = 16'b11111_101110_00000;
    timing1[2][12] = 16'b00000_000000_00000;
    timing1[2][13] = 16'b00000_000000_00000;
    timing1[2][14] = 16'b11111_111110_11111;
    timing1[3][0] = 16'b11111_111110_11111;
    timing1[3][1] = 16'b00000_000000_00000;
    timing1[3][2] = 16'b11111_101110_00000;
    timing1[3][3] = 16'b11111_101110_00000;
    timing1[3][4] = 16'b11001_100100_00000;
    timing1[3][5] = 16'b11111_111110_11111;
    timing1[3][6] = 16'b11111_111110_11111;
    timing1[3][7] = 16'b00111_001111_00111;
    timing1[3][8] = 16'b11111_111110_11111;
    timing1[3][9] = 16'b11111_111110_11111;
    timing1[3][10] = 16'b11001_100100_00000;
    timing1[3][11] = 16'b11111_101110_00000;
    timing1[3][12] = 16'b11111_101110_00000;
    timing1[3][13] = 16'b00000_000000_00000;
    timing1[3][14] = 16'b11111_111110_11111;
    timing1[4][0] = 16'b11111_111110_11111;
    timing1[4][1] = 16'b00000_000000_00000;
    timing1[4][2] = 16'b11111_101110_00000;
    timing1[4][3] = 16'b11001_100100_00000;
    timing1[4][4] = 16'b11111_111110_11111;
    timing1[4][5] = 16'b11111_111110_11111;
    timing1[4][6] = 16'b11111_111110_11111;
    timing1[4][7] = 16'b00111_001111_00111;
    timing1[4][8] = 16'b11111_111110_11111;
    timing1[4][9] = 16'b11111_111110_11111;
    timing1[4][10] = 16'b11111_111110_11111;
    timing1[4][11] = 16'b11001_100100_00000;
    timing1[4][12] = 16'b11111_101110_00000;
    timing1[4][13] = 16'b00000_000000_00000;
    timing1[4][14] = 16'b11111_111110_11111;
    timing1[5][0] = 16'b11111_111110_11111;
    timing1[5][1] = 16'b11111_101110_00000;
    timing1[5][2] = 16'b11001_100100_00000;
    timing1[5][3] = 16'b11111_111110_11111;
    timing1[5][4] = 16'b11111_111110_11111;
    timing1[5][5] = 16'b11111_111110_11111;
    timing1[5][6] = 16'b11111_111110_11111;
    timing1[5][7] = 16'b00111_001111_00111;
    timing1[5][8] = 16'b11111_111110_11111;
    timing1[5][9] = 16'b11111_111110_11111;
    timing1[5][10] = 16'b11111_111110_11111;
    timing1[5][11] = 16'b11111_111110_11111;
    timing1[5][12] = 16'b11001_100100_00000;
    timing1[5][13] = 16'b11111_101110_00000;
    timing1[5][14] = 16'b11111_111110_11111;
    timing1[6][0] = 16'b11111_111110_11111;
    timing1[6][1] = 16'b11111_101110_00000;
    timing1[6][2] = 16'b11001_100100_00000;
    timing1[6][3] = 16'b11111_111110_11111;
    timing1[6][4] = 16'b11111_111110_11111;
    timing1[6][5] = 16'b11111_111110_11111;
    timing1[6][6] = 16'b11111_111110_11111;
    timing1[6][7] = 16'b00111_001111_00111;
    timing1[6][8] = 16'b11111_111110_11111;
    timing1[6][9] = 16'b11111_111110_11111;
    timing1[6][10] = 16'b11111_111110_11111;
    timing1[6][11] = 16'b11111_111110_11111;
    timing1[6][12] = 16'b11001_100100_00000;
    timing1[6][13] = 16'b11111_101110_00000;
    timing1[6][14] = 16'b11111_111110_11111;
    timing1[7][0] = 16'b11111_111110_11111;
    timing1[7][1] = 16'b11111_101110_00000;
    timing1[7][2] = 16'b11001_100100_00000;
    timing1[7][3] = 16'b11111_111110_11111;
    timing1[7][4] = 16'b11111_111110_11111;
    timing1[7][5] = 16'b11111_111110_11111;
    timing1[7][6] = 16'b11111_111110_11111;
    timing1[7][7] = 16'b00000_000000_00000;
    timing1[7][8] = 16'b00000_000000_00000;
    timing1[7][9] = 16'b00000_000000_00000;
    timing1[7][10] = 16'b00000_000000_00000;
    timing1[7][11] = 16'b11111_111110_11111;
    timing1[7][12] = 16'b11001_100100_00000;
    timing1[7][13] = 16'b11111_101110_00000;
    timing1[7][14] = 16'b11111_111110_11111;
    timing1[8][0] = 16'b11111_111110_11111;
    timing1[8][1] = 16'b11111_101110_00000;
    timing1[8][2] = 16'b11001_100100_00000;
    timing1[8][3] = 16'b11111_111110_11111;
    timing1[8][4] = 16'b11111_111110_11111;
    timing1[8][5] = 16'b11111_111110_11111;
    timing1[8][6] = 16'b11111_111110_11111;
    timing1[8][7] = 16'b11111_111110_11111;
    timing1[8][8] = 16'b11111_111110_11111;
    timing1[8][9] = 16'b11111_111110_11111;
    timing1[8][10] = 16'b11111_111110_11111;
    timing1[8][11] = 16'b11111_111110_11111;
    timing1[8][12] = 16'b11001_100100_00000;
    timing1[8][13] = 16'b11111_101110_00000;
    timing1[8][14] = 16'b11111_111110_11111;
    timing1[9][0] = 16'b11111_111110_11111;
    timing1[9][1] = 16'b11111_101110_00000;
    timing1[9][2] = 16'b11001_100100_00000;
    timing1[9][3] = 16'b11111_111110_11111;
    timing1[9][4] = 16'b11111_111110_11111;
    timing1[9][5] = 16'b11111_111110_11111;
    timing1[9][6] = 16'b11111_111110_11111;
    timing1[9][7] = 16'b11111_111110_11111;
    timing1[9][8] = 16'b11111_111110_11111;
    timing1[9][9] = 16'b11111_111110_11111;
    timing1[9][10] = 16'b11111_111110_11111;
    timing1[9][11] = 16'b11111_111110_11111;
    timing1[9][12] = 16'b11001_100100_00000;
    timing1[9][13] = 16'b11111_101110_00000;
    timing1[9][14] = 16'b11111_111110_11111;
    timing1[10][0] = 16'b11111_111110_11111;
    timing1[10][1] = 16'b00000_000000_00000;
    timing1[10][2] = 16'b11111_101110_00000;
    timing1[10][3] = 16'b11001_100100_00000;
    timing1[10][4] = 16'b11111_111110_11111;
    timing1[10][5] = 16'b11111_111110_11111;
    timing1[10][6] = 16'b11111_111110_11111;
    timing1[10][7] = 16'b11111_111110_11111;
    timing1[10][8] = 16'b11111_111110_11111;
    timing1[10][9] = 16'b11111_111110_11111;
    timing1[10][10] = 16'b11111_111110_11111;
    timing1[10][11] = 16'b11001_100100_00000;
    timing1[10][12] = 16'b11111_101110_00000;
    timing1[10][13] = 16'b00000_000000_00000;
    timing1[10][14] = 16'b11111_111110_11111;
    timing1[11][0] = 16'b11111_111110_11111;
    timing1[11][1] = 16'b00000_000000_00000;
    timing1[11][2] = 16'b11111_101110_00000;
    timing1[11][3] = 16'b11111_101110_00000;
    timing1[11][4] = 16'b11001_100100_00000;
    timing1[11][5] = 16'b11111_111110_11111;
    timing1[11][6] = 16'b11111_111110_11111;
    timing1[11][7] = 16'b11111_111110_11111;
    timing1[11][8] = 16'b11111_111110_11111;
    timing1[11][9] = 16'b11111_111110_11111;
    timing1[11][10] = 16'b11001_100100_00000;
    timing1[11][11] = 16'b11111_101110_00000;
    timing1[11][12] = 16'b11111_101110_00000;
    timing1[11][13] = 16'b00000_000000_00000;
    timing1[11][14] = 16'b11111_111110_11111;
    timing1[12][0] = 16'b11111_111110_11111;
    timing1[12][1] = 16'b00000_000000_00000;
    timing1[12][2] = 16'b00000_000000_00000;
    timing1[12][3] = 16'b11111_101110_00000;
    timing1[12][4] = 16'b11111_101110_00000;
    timing1[12][5] = 16'b11001_100100_00000;
    timing1[12][6] = 16'b11001_100100_00000;
    timing1[12][7] = 16'b11001_100100_00000;
    timing1[12][8] = 16'b11001_100100_00000;
    timing1[12][9] = 16'b11001_100100_00000;
    timing1[12][10] = 16'b11111_101110_00000;
    timing1[12][11] = 16'b11111_101110_00000;
    timing1[12][12] = 16'b00000_000000_00000;
    timing1[12][13] = 16'b00000_000000_00000;
    timing1[12][14] = 16'b11111_111110_11111;
    timing1[13][0] = 16'b11111_111110_11111;
    timing1[13][1] = 16'b00000_000000_00000;
    timing1[13][2] = 16'b00000_000000_00000;
    timing1[13][3] = 16'b00000_000000_00000;
    timing1[13][4] = 16'b00000_000000_00000;
    timing1[13][5] = 16'b11111_101110_00000;
    timing1[13][6] = 16'b11111_101110_00000;
    timing1[13][7] = 16'b11111_101110_00000;
    timing1[13][8] = 16'b11111_101110_00000;
    timing1[13][9] = 16'b11111_101110_00000;
    timing1[13][10] = 16'b00000_000000_00000;
    timing1[13][11] = 16'b00000_000000_00000;
    timing1[13][12] = 16'b00000_000000_00000;
    timing1[13][13] = 16'b00000_000000_00000;
    timing1[13][14] = 16'b11111_111110_11111;
    timing1[14][0] = 16'b11111_111110_11111;
    timing1[14][1] = 16'b11111_111110_11111;
    timing1[14][2] = 16'b11111_111110_11111;
    timing1[14][3] = 16'b11111_111110_11111;
    timing1[14][4] = 16'b11111_111110_11111;
    timing1[14][5] = 16'b11111_111110_11111;
    timing1[14][6] = 16'b11111_111110_11111;
    timing1[14][7] = 16'b11111_111110_11111;
    timing1[14][8] = 16'b11111_111110_11111;
    timing1[14][9] = 16'b11111_111110_11111;
    timing1[14][10] = 16'b11111_111110_11111;
    timing1[14][11] = 16'b11111_111110_11111;
    timing1[14][12] = 16'b11111_111110_11111;
    timing1[14][13] = 16'b11111_111110_11111;
    timing1[14][14] = 16'b11111_111110_11111;
    
    timing2[0][0] = 16'b11111_111110_11111;
    timing2[0][1] = 16'b11111_111110_11111;
    timing2[0][2] = 16'b11111_111110_11111;
    timing2[0][3] = 16'b11111_111110_11111;
    timing2[0][4] = 16'b11111_111110_11111;
    timing2[0][5] = 16'b11111_111110_11111;
    timing2[0][6] = 16'b11111_111110_11111;
    timing2[0][7] = 16'b11111_111110_11111;
    timing2[0][8] = 16'b11111_111110_11111;
    timing2[0][9] = 16'b11111_111110_11111;
    timing2[0][10] = 16'b11111_111110_11111;
    timing2[0][11] = 16'b11111_111110_11111;
    timing2[0][12] = 16'b11111_111110_11111;
    timing2[0][13] = 16'b11111_111110_11111;
    timing2[0][14] = 16'b11111_111110_11111;
    timing2[1][0] = 16'b11111_111110_11111;
    timing2[1][1] = 16'b00000_000000_00000;
    timing2[1][2] = 16'b00000_000000_00000;
    timing2[1][3] = 16'b00000_000000_00000;
    timing2[1][4] = 16'b00000_000000_00000;
    timing2[1][5] = 16'b11111_101110_00000;
    timing2[1][6] = 16'b11111_101110_00000;
    timing2[1][7] = 16'b11111_101110_00000;
    timing2[1][8] = 16'b11111_101110_00000;
    timing2[1][9] = 16'b11111_101110_00000;
    timing2[1][10] = 16'b00000_000000_00000;
    timing2[1][11] = 16'b00000_000000_00000;
    timing2[1][12] = 16'b00000_000000_00000;
    timing2[1][13] = 16'b00000_000000_00000;
    timing2[1][14] = 16'b11111_111110_11111;
    timing2[2][0] = 16'b11111_111110_11111;
    timing2[2][1] = 16'b00000_000000_00000;
    timing2[2][2] = 16'b00000_000000_00000;
    timing2[2][3] = 16'b11111_101110_00000;
    timing2[2][4] = 16'b11111_101110_00000;
    timing2[2][5] = 16'b11001_100100_00000;
    timing2[2][6] = 16'b11001_100100_00000;
    timing2[2][7] = 16'b11001_100100_00000;
    timing2[2][8] = 16'b11001_100100_00000;
    timing2[2][9] = 16'b11001_100100_00000;
    timing2[2][10] = 16'b11111_101110_00000;
    timing2[2][11] = 16'b11111_101110_00000;
    timing2[2][12] = 16'b00000_000000_00000;
    timing2[2][13] = 16'b00000_000000_00000;
    timing2[2][14] = 16'b11111_111110_11111;
    timing2[3][0] = 16'b11111_111110_11111;
    timing2[3][1] = 16'b00000_000000_00000;
    timing2[3][2] = 16'b11111_101110_00000;
    timing2[3][3] = 16'b11111_101110_00000;
    timing2[3][4] = 16'b11001_100100_00000;
    timing2[3][5] = 16'b11111_111110_11111;
    timing2[3][6] = 16'b11111_111110_11111;
    timing2[3][7] = 16'b11111_111110_11111;
    timing2[3][8] = 16'b11111_111110_11111;
    timing2[3][9] = 16'b11111_111110_11111;
    timing2[3][10] = 16'b11001_100100_00000;
    timing2[3][11] = 16'b11111_101110_00000;
    timing2[3][12] = 16'b11111_101110_00000;
    timing2[3][13] = 16'b00000_000000_00000;
    timing2[3][14] = 16'b11111_111110_11111;
    timing2[4][0] = 16'b11111_111110_11111;
    timing2[4][1] = 16'b00000_000000_00000;
    timing2[4][2] = 16'b11111_101110_00000;
    timing2[4][3] = 16'b11001_100100_00000;
    timing2[4][4] = 16'b11111_111110_11111;
    timing2[4][5] = 16'b11111_111110_11111;
    timing2[4][6] = 16'b11111_111110_11111;
    timing2[4][7] = 16'b11111_111110_11111;
    timing2[4][8] = 16'b11111_111110_11111;
    timing2[4][9] = 16'b00111_001111_00111;
    timing2[4][10] = 16'b11111_111110_11111;
    timing2[4][11] = 16'b11001_100100_00000;
    timing2[4][12] = 16'b11111_101110_00000;
    timing2[4][13] = 16'b00000_000000_00000;
    timing2[4][14] = 16'b11111_111110_11111;
    timing2[5][0] = 16'b11111_111110_11111;
    timing2[5][1] = 16'b11111_101110_00000;
    timing2[5][2] = 16'b11001_100100_00000;
    timing2[5][3] = 16'b11111_111110_11111;
    timing2[5][4] = 16'b11111_111110_11111;
    timing2[5][5] = 16'b11111_111110_11111;
    timing2[5][6] = 16'b11111_111110_11111;
    timing2[5][7] = 16'b11111_111110_11111;
    timing2[5][8] = 16'b11111_111110_11111;
    timing2[5][9] = 16'b00111_001111_00111;
    timing2[5][10] = 16'b11111_111110_11111;
    timing2[5][11] = 16'b11111_111110_11111;
    timing2[5][12] = 16'b11001_100100_00000;
    timing2[5][13] = 16'b11111_101110_00000;
    timing2[5][14] = 16'b11111_111110_11111;
    timing2[6][0] = 16'b11111_111110_11111;
    timing2[6][1] = 16'b11111_101110_00000;
    timing2[6][2] = 16'b11001_100100_00000;
    timing2[6][3] = 16'b11111_111110_11111;
    timing2[6][4] = 16'b11111_111110_11111;
    timing2[6][5] = 16'b11111_111110_11111;
    timing2[6][6] = 16'b11111_111110_11111;
    timing2[6][7] = 16'b11111_111110_11111;
    timing2[6][8] = 16'b00111_001111_00111;
    timing2[6][9] = 16'b11111_111110_11111;
    timing2[6][10] = 16'b11111_111110_11111;
    timing2[6][11] = 16'b11111_111110_11111;
    timing2[6][12] = 16'b11001_100100_00000;
    timing2[6][13] = 16'b11111_101110_00000;
    timing2[6][14] = 16'b11111_111110_11111;
    timing2[7][0] = 16'b11111_111110_11111;
    timing2[7][1] = 16'b11111_101110_00000;
    timing2[7][2] = 16'b11001_100100_00000;
    timing2[7][3] = 16'b11111_111110_11111;
    timing2[7][4] = 16'b11111_111110_11111;
    timing2[7][5] = 16'b11111_111110_11111;
    timing2[7][6] = 16'b11111_111110_11111;
    timing2[7][7] = 16'b00000_000000_00000;
    timing2[7][8] = 16'b00000_000000_00000;
    timing2[7][9] = 16'b00000_000000_00000;
    timing2[7][10] = 16'b00000_000000_00000;
    timing2[7][11] = 16'b11111_111110_11111;
    timing2[7][12] = 16'b11001_100100_00000;
    timing2[7][13] = 16'b11111_101110_00000;
    timing2[7][14] = 16'b11111_111110_11111;
    timing2[8][0] = 16'b11111_111110_11111;
    timing2[8][1] = 16'b11111_101110_00000;
    timing2[8][2] = 16'b11001_100100_00000;
    timing2[8][3] = 16'b11111_111110_11111;
    timing2[8][4] = 16'b11111_111110_11111;
    timing2[8][5] = 16'b11111_111110_11111;
    timing2[8][6] = 16'b11111_111110_11111;
    timing2[8][7] = 16'b11111_111110_11111;
    timing2[8][8] = 16'b11111_111110_11111;
    timing2[8][9] = 16'b11111_111110_11111;
    timing2[8][10] = 16'b11111_111110_11111;
    timing2[8][11] = 16'b11111_111110_11111;
    timing2[8][12] = 16'b11001_100100_00000;
    timing2[8][13] = 16'b11111_101110_00000;
    timing2[8][14] = 16'b11111_111110_11111;
    timing2[9][0] = 16'b11111_111110_11111;
    timing2[9][1] = 16'b11111_101110_00000;
    timing2[9][2] = 16'b11001_100100_00000;
    timing2[9][3] = 16'b11111_111110_11111;
    timing2[9][4] = 16'b11111_111110_11111;
    timing2[9][5] = 16'b11111_111110_11111;
    timing2[9][6] = 16'b11111_111110_11111;
    timing2[9][7] = 16'b11111_111110_11111;
    timing2[9][8] = 16'b11111_111110_11111;
    timing2[9][9] = 16'b11111_111110_11111;
    timing2[9][10] = 16'b11111_111110_11111;
    timing2[9][11] = 16'b11111_111110_11111;
    timing2[9][12] = 16'b11001_100100_00000;
    timing2[9][13] = 16'b11111_101110_00000;
    timing2[9][14] = 16'b11111_111110_11111;
    timing2[10][0] = 16'b11111_111110_11111;
    timing2[10][1] = 16'b00000_000000_00000;
    timing2[10][2] = 16'b11111_101110_00000;
    timing2[10][3] = 16'b11001_100100_00000;
    timing2[10][4] = 16'b11111_111110_11111;
    timing2[10][5] = 16'b11111_111110_11111;
    timing2[10][6] = 16'b11111_111110_11111;
    timing2[10][7] = 16'b11111_111110_11111;
    timing2[10][8] = 16'b11111_111110_11111;
    timing2[10][9] = 16'b11111_111110_11111;
    timing2[10][10] = 16'b11111_111110_11111;
    timing2[10][11] = 16'b11001_100100_00000;
    timing2[10][12] = 16'b11111_101110_00000;
    timing2[10][13] = 16'b00000_000000_00000;
    timing2[10][14] = 16'b11111_111110_11111;
    timing2[11][0] = 16'b11111_111110_11111;
    timing2[11][1] = 16'b00000_000000_00000;
    timing2[11][2] = 16'b11111_101110_00000;
    timing2[11][3] = 16'b11111_101110_00000;
    timing2[11][4] = 16'b11001_100100_00000;
    timing2[11][5] = 16'b11111_111110_11111;
    timing2[11][6] = 16'b11111_111110_11111;
    timing2[11][7] = 16'b11111_111110_11111;
    timing2[11][8] = 16'b11111_111110_11111;
    timing2[11][9] = 16'b11111_111110_11111;
    timing2[11][10] = 16'b11001_100100_00000;
    timing2[11][11] = 16'b11111_101110_00000;
    timing2[11][12] = 16'b11111_101110_00000;
    timing2[11][13] = 16'b00000_000000_00000;
    timing2[11][14] = 16'b11111_111110_11111;
    timing2[12][0] = 16'b11111_111110_11111;
    timing2[12][1] = 16'b00000_000000_00000;
    timing2[12][2] = 16'b00000_000000_00000;
    timing2[12][3] = 16'b11111_101110_00000;
    timing2[12][4] = 16'b11111_101110_00000;
    timing2[12][5] = 16'b11001_100100_00000;
    timing2[12][6] = 16'b11001_100100_00000;
    timing2[12][7] = 16'b11001_100100_00000;
    timing2[12][8] = 16'b11001_100100_00000;
    timing2[12][9] = 16'b11001_100100_00000;
    timing2[12][10] = 16'b11111_101110_00000;
    timing2[12][11] = 16'b11111_101110_00000;
    timing2[12][12] = 16'b00000_000000_00000;
    timing2[12][13] = 16'b00000_000000_00000;
    timing2[12][14] = 16'b11111_111110_11111;
    timing2[13][0] = 16'b11111_111110_11111;
    timing2[13][1] = 16'b00000_000000_00000;
    timing2[13][2] = 16'b00000_000000_00000;
    timing2[13][3] = 16'b00000_000000_00000;
    timing2[13][4] = 16'b00000_000000_00000;
    timing2[13][5] = 16'b11111_101110_00000;
    timing2[13][6] = 16'b11111_101110_00000;
    timing2[13][7] = 16'b11111_101110_00000;
    timing2[13][8] = 16'b11111_101110_00000;
    timing2[13][9] = 16'b11111_101110_00000;
    timing2[13][10] = 16'b00000_000000_00000;
    timing2[13][11] = 16'b00000_000000_00000;
    timing2[13][12] = 16'b00000_000000_00000;
    timing2[13][13] = 16'b00000_000000_00000;
    timing2[13][14] = 16'b11111_111110_11111;
    timing2[14][0] = 16'b11111_111110_11111;
    timing2[14][1] = 16'b11111_111110_11111;
    timing2[14][2] = 16'b11111_111110_11111;
    timing2[14][3] = 16'b11111_111110_11111;
    timing2[14][4] = 16'b11111_111110_11111;
    timing2[14][5] = 16'b11111_111110_11111;
    timing2[14][6] = 16'b11111_111110_11111;
    timing2[14][7] = 16'b11111_111110_11111;
    timing2[14][8] = 16'b11111_111110_11111;
    timing2[14][9] = 16'b11111_111110_11111;
    timing2[14][10] = 16'b11111_111110_11111;
    timing2[14][11] = 16'b11111_111110_11111;
    timing2[14][12] = 16'b11111_111110_11111;
    timing2[14][13] = 16'b11111_111110_11111;
    timing2[14][14] = 16'b11111_111110_11111;
    
    timing3[0][0] = 16'b11111_111110_11111;
    timing3[0][1] = 16'b11111_111110_11111;
    timing3[0][2] = 16'b11111_111110_11111;
    timing3[0][3] = 16'b11111_111110_11111;
    timing3[0][4] = 16'b11111_111110_11111;
    timing3[0][5] = 16'b11111_111110_11111;
    timing3[0][6] = 16'b11111_111110_11111;
    timing3[0][7] = 16'b11111_111110_11111;
    timing3[0][8] = 16'b11111_111110_11111;
    timing3[0][9] = 16'b11111_111110_11111;
    timing3[0][10] = 16'b11111_111110_11111;
    timing3[0][11] = 16'b11111_111110_11111;
    timing3[0][12] = 16'b11111_111110_11111;
    timing3[0][13] = 16'b11111_111110_11111;
    timing3[0][14] = 16'b11111_111110_11111;
    timing3[1][0] = 16'b11111_111110_11111;
    timing3[1][1] = 16'b00000_000000_00000;
    timing3[1][2] = 16'b00000_000000_00000;
    timing3[1][3] = 16'b00000_000000_00000;
    timing3[1][4] = 16'b00000_000000_00000;
    timing3[1][5] = 16'b11111_101110_00000;
    timing3[1][6] = 16'b11111_101110_00000;
    timing3[1][7] = 16'b11111_101110_00000;
    timing3[1][8] = 16'b11111_101110_00000;
    timing3[1][9] = 16'b11111_101110_00000;
    timing3[1][10] = 16'b00000_000000_00000;
    timing3[1][11] = 16'b00000_000000_00000;
    timing3[1][12] = 16'b00000_000000_00000;
    timing3[1][13] = 16'b00000_000000_00000;
    timing3[1][14] = 16'b11111_111110_11111;
    timing3[2][0] = 16'b11111_111110_11111;
    timing3[2][1] = 16'b00000_000000_00000;
    timing3[2][2] = 16'b00000_000000_00000;
    timing3[2][3] = 16'b11111_101110_00000;
    timing3[2][4] = 16'b11111_101110_00000;
    timing3[2][5] = 16'b11001_100100_00000;
    timing3[2][6] = 16'b11001_100100_00000;
    timing3[2][7] = 16'b11001_100100_00000;
    timing3[2][8] = 16'b11001_100100_00000;
    timing3[2][9] = 16'b11001_100100_00000;
    timing3[2][10] = 16'b11111_101110_00000;
    timing3[2][11] = 16'b11111_101110_00000;
    timing3[2][12] = 16'b00000_000000_00000;
    timing3[2][13] = 16'b00000_000000_00000;
    timing3[2][14] = 16'b11111_111110_11111;
    timing3[3][0] = 16'b11111_111110_11111;
    timing3[3][1] = 16'b00000_000000_00000;
    timing3[3][2] = 16'b11111_101110_00000;
    timing3[3][3] = 16'b11111_101110_00000;
    timing3[3][4] = 16'b11001_100100_00000;
    timing3[3][5] = 16'b11111_111110_11111;
    timing3[3][6] = 16'b11111_111110_11111;
    timing3[3][7] = 16'b11111_111110_11111;
    timing3[3][8] = 16'b11111_111110_11111;
    timing3[3][9] = 16'b11111_111110_11111;
    timing3[3][10] = 16'b11001_100100_00000;
    timing3[3][11] = 16'b11111_101110_00000;
    timing3[3][12] = 16'b11111_101110_00000;
    timing3[3][13] = 16'b00000_000000_00000;
    timing3[3][14] = 16'b11111_111110_11111;
    timing3[4][0] = 16'b11111_111110_11111;
    timing3[4][1] = 16'b00000_000000_00000;
    timing3[4][2] = 16'b11111_101110_00000;
    timing3[4][3] = 16'b11001_100100_00000;
    timing3[4][4] = 16'b11111_111110_11111;
    timing3[4][5] = 16'b11111_111110_11111;
    timing3[4][6] = 16'b11111_111110_11111;
    timing3[4][7] = 16'b11111_111110_11111;
    timing3[4][8] = 16'b11111_111110_11111;
    timing3[4][9] = 16'b11111_111110_11111;
    timing3[4][10] = 16'b11111_111110_11111;
    timing3[4][11] = 16'b11001_100100_00000;
    timing3[4][12] = 16'b11111_101110_00000;
    timing3[4][13] = 16'b00000_000000_00000;
    timing3[4][14] = 16'b11111_111110_11111;
    timing3[5][0] = 16'b11111_111110_11111;
    timing3[5][1] = 16'b11111_101110_00000;
    timing3[5][2] = 16'b11001_100100_00000;
    timing3[5][3] = 16'b11111_111110_11111;
    timing3[5][4] = 16'b11111_111110_11111;
    timing3[5][5] = 16'b11111_111110_11111;
    timing3[5][6] = 16'b11111_111110_11111;
    timing3[5][7] = 16'b11111_111110_11111;
    timing3[5][8] = 16'b11111_111110_11111;
    timing3[5][9] = 16'b11111_111110_11111;
    timing3[5][10] = 16'b11111_111110_11111;
    timing3[5][11] = 16'b11111_111110_11111;
    timing3[5][12] = 16'b11001_100100_00000;
    timing3[5][13] = 16'b11111_101110_00000;
    timing3[5][14] = 16'b11111_111110_11111;
    timing3[6][0] = 16'b11111_111110_11111;
    timing3[6][1] = 16'b11111_101110_00000;
    timing3[6][2] = 16'b11001_100100_00000;
    timing3[6][3] = 16'b11111_111110_11111;
    timing3[6][4] = 16'b11111_111110_11111;
    timing3[6][5] = 16'b11111_111110_11111;
    timing3[6][6] = 16'b11111_111110_11111;
    timing3[6][7] = 16'b11111_111110_11111;
    timing3[6][8] = 16'b11111_111110_11111;
    timing3[6][9] = 16'b11111_111110_11111;
    timing3[6][10] = 16'b11111_111110_11111;
    timing3[6][11] = 16'b11111_111110_11111;
    timing3[6][12] = 16'b11001_100100_00000;
    timing3[6][13] = 16'b11111_101110_00000;
    timing3[6][14] = 16'b11111_111110_11111;
    timing3[7][0] = 16'b11111_111110_11111;
    timing3[7][1] = 16'b11111_101110_00000;
    timing3[7][2] = 16'b11001_100100_00000;
    timing3[7][3] = 16'b11111_111110_11111;
    timing3[7][4] = 16'b11111_111110_11111;
    timing3[7][5] = 16'b11111_111110_11111;
    timing3[7][6] = 16'b11111_111110_11111;
    timing3[7][7] = 16'b00000_000000_00000;
    timing3[7][8] = 16'b00000_000000_00000;
    timing3[7][9] = 16'b00000_000000_00000;
    timing3[7][10] = 16'b00000_000000_00000;
    timing3[7][11] = 16'b00111_001111_00111;
    timing3[7][12] = 16'b11001_100100_00000;
    timing3[7][13] = 16'b11111_101110_00000;
    timing3[7][14] = 16'b11111_111110_11111;
    timing3[8][0] = 16'b11111_111110_11111;
    timing3[8][1] = 16'b11111_101110_00000;
    timing3[8][2] = 16'b11001_100100_00000;
    timing3[8][3] = 16'b11111_111110_11111;
    timing3[8][4] = 16'b11111_111110_11111;
    timing3[8][5] = 16'b11111_111110_11111;
    timing3[8][6] = 16'b11111_111110_11111;
    timing3[8][7] = 16'b11111_111110_11111;
    timing3[8][8] = 16'b11111_111110_11111;
    timing3[8][9] = 16'b11111_111110_11111;
    timing3[8][10] = 16'b11111_111110_11111;
    timing3[8][11] = 16'b11111_111110_11111;
    timing3[8][12] = 16'b11001_100100_00000;
    timing3[8][13] = 16'b11111_101110_00000;
    timing3[8][14] = 16'b11111_111110_11111;
    timing3[9][0] = 16'b11111_111110_11111;
    timing3[9][1] = 16'b11111_101110_00000;
    timing3[9][2] = 16'b11001_100100_00000;
    timing3[9][3] = 16'b11111_111110_11111;
    timing3[9][4] = 16'b11111_111110_11111;
    timing3[9][5] = 16'b11111_111110_11111;
    timing3[9][6] = 16'b11111_111110_11111;
    timing3[9][7] = 16'b11111_111110_11111;
    timing3[9][8] = 16'b11111_111110_11111;
    timing3[9][9] = 16'b11111_111110_11111;
    timing3[9][10] = 16'b11111_111110_11111;
    timing3[9][11] = 16'b11111_111110_11111;
    timing3[9][12] = 16'b11001_100100_00000;
    timing3[9][13] = 16'b11111_101110_00000;
    timing3[9][14] = 16'b11111_111110_11111;
    timing3[10][0] = 16'b11111_111110_11111;
    timing3[10][1] = 16'b00000_000000_00000;
    timing3[10][2] = 16'b11111_101110_00000;
    timing3[10][3] = 16'b11001_100100_00000;
    timing3[10][4] = 16'b11111_111110_11111;
    timing3[10][5] = 16'b11111_111110_11111;
    timing3[10][6] = 16'b11111_111110_11111;
    timing3[10][7] = 16'b11111_111110_11111;
    timing3[10][8] = 16'b11111_111110_11111;
    timing3[10][9] = 16'b11111_111110_11111;
    timing3[10][10] = 16'b11111_111110_11111;
    timing3[10][11] = 16'b11001_100100_00000;
    timing3[10][12] = 16'b11111_101110_00000;
    timing3[10][13] = 16'b00000_000000_00000;
    timing3[10][14] = 16'b11111_111110_11111;
    timing3[11][0] = 16'b11111_111110_11111;
    timing3[11][1] = 16'b00000_000000_00000;
    timing3[11][2] = 16'b11111_101110_00000;
    timing3[11][3] = 16'b11111_101110_00000;
    timing3[11][4] = 16'b11001_100100_00000;
    timing3[11][5] = 16'b11111_111110_11111;
    timing3[11][6] = 16'b11111_111110_11111;
    timing3[11][7] = 16'b11111_111110_11111;
    timing3[11][8] = 16'b11111_111110_11111;
    timing3[11][9] = 16'b11111_111110_11111;
    timing3[11][10] = 16'b11001_100100_00000;
    timing3[11][11] = 16'b11111_101110_00000;
    timing3[11][12] = 16'b11111_101110_00000;
    timing3[11][13] = 16'b00000_000000_00000;
    timing3[11][14] = 16'b11111_111110_11111;
    timing3[12][0] = 16'b11111_111110_11111;
    timing3[12][1] = 16'b00000_000000_00000;
    timing3[12][2] = 16'b00000_000000_00000;
    timing3[12][3] = 16'b11111_101110_00000;
    timing3[12][4] = 16'b11111_101110_00000;
    timing3[12][5] = 16'b11001_100100_00000;
    timing3[12][6] = 16'b11001_100100_00000;
    timing3[12][7] = 16'b11001_100100_00000;
    timing3[12][8] = 16'b11001_100100_00000;
    timing3[12][9] = 16'b11001_100100_00000;
    timing3[12][10] = 16'b11111_101110_00000;
    timing3[12][11] = 16'b11111_101110_00000;
    timing3[12][12] = 16'b00000_000000_00000;
    timing3[12][13] = 16'b00000_000000_00000;
    timing3[12][14] = 16'b11111_111110_11111;
    timing3[13][0] = 16'b11111_111110_11111;
    timing3[13][1] = 16'b00000_000000_00000;
    timing3[13][2] = 16'b00000_000000_00000;
    timing3[13][3] = 16'b00000_000000_00000;
    timing3[13][4] = 16'b00000_000000_00000;
    timing3[13][5] = 16'b11111_101110_00000;
    timing3[13][6] = 16'b11111_101110_00000;
    timing3[13][7] = 16'b11111_101110_00000;
    timing3[13][8] = 16'b11111_101110_00000;
    timing3[13][9] = 16'b11111_101110_00000;
    timing3[13][10] = 16'b00000_000000_00000;
    timing3[13][11] = 16'b00000_000000_00000;
    timing3[13][12] = 16'b00000_000000_00000;
    timing3[13][13] = 16'b00000_000000_00000;
    timing3[13][14] = 16'b11111_111110_11111;
    timing3[14][0] = 16'b11111_111110_11111;
    timing3[14][1] = 16'b11111_111110_11111;
    timing3[14][2] = 16'b11111_111110_11111;
    timing3[14][3] = 16'b11111_111110_11111;
    timing3[14][4] = 16'b11111_111110_11111;
    timing3[14][5] = 16'b11111_111110_11111;
    timing3[14][6] = 16'b11111_111110_11111;
    timing3[14][7] = 16'b11111_111110_11111;
    timing3[14][8] = 16'b11111_111110_11111;
    timing3[14][9] = 16'b11111_111110_11111;
    timing3[14][10] = 16'b11111_111110_11111;
    timing3[14][11] = 16'b11111_111110_11111;
    timing3[14][12] = 16'b11111_111110_11111;
    timing3[14][13] = 16'b11111_111110_11111;
    timing3[14][14] = 16'b11111_111110_11111;
    
    timing4[0][0] = 16'b11111_111110_11111;
    timing4[0][1] = 16'b11111_111110_11111;
    timing4[0][2] = 16'b11111_111110_11111;
    timing4[0][3] = 16'b11111_111110_11111;
    timing4[0][4] = 16'b11111_111110_11111;
    timing4[0][5] = 16'b11111_111110_11111;
    timing4[0][6] = 16'b11111_111110_11111;
    timing4[0][7] = 16'b11111_111110_11111;
    timing4[0][8] = 16'b11111_111110_11111;
    timing4[0][9] = 16'b11111_111110_11111;
    timing4[0][10] = 16'b11111_111110_11111;
    timing4[0][11] = 16'b11111_111110_11111;
    timing4[0][12] = 16'b11111_111110_11111;
    timing4[0][13] = 16'b11111_111110_11111;
    timing4[0][14] = 16'b11111_111110_11111;
    timing4[1][0] = 16'b11111_111110_11111;
    timing4[1][1] = 16'b00000_000000_00000;
    timing4[1][2] = 16'b00000_000000_00000;
    timing4[1][3] = 16'b00000_000000_00000;
    timing4[1][4] = 16'b00000_000000_00000;
    timing4[1][5] = 16'b11111_101110_00000;
    timing4[1][6] = 16'b11111_101110_00000;
    timing4[1][7] = 16'b11111_101110_00000;
    timing4[1][8] = 16'b11111_101110_00000;
    timing4[1][9] = 16'b11111_101110_00000;
    timing4[1][10] = 16'b00000_000000_00000;
    timing4[1][11] = 16'b00000_000000_00000;
    timing4[1][12] = 16'b00000_000000_00000;
    timing4[1][13] = 16'b00000_000000_00000;
    timing4[1][14] = 16'b11111_111110_11111;
    timing4[2][0] = 16'b11111_111110_11111;
    timing4[2][1] = 16'b00000_000000_00000;
    timing4[2][2] = 16'b00000_000000_00000;
    timing4[2][3] = 16'b11111_101110_00000;
    timing4[2][4] = 16'b11111_101110_00000;
    timing4[2][5] = 16'b11001_100100_00000;
    timing4[2][6] = 16'b11001_100100_00000;
    timing4[2][7] = 16'b11001_100100_00000;
    timing4[2][8] = 16'b11001_100100_00000;
    timing4[2][9] = 16'b11001_100100_00000;
    timing4[2][10] = 16'b11111_101110_00000;
    timing4[2][11] = 16'b11111_101110_00000;
    timing4[2][12] = 16'b00000_000000_00000;
    timing4[2][13] = 16'b00000_000000_00000;
    timing4[2][14] = 16'b11111_111110_11111;
    timing4[3][0] = 16'b11111_111110_11111;
    timing4[3][1] = 16'b00000_000000_00000;
    timing4[3][2] = 16'b11111_101110_00000;
    timing4[3][3] = 16'b11111_101110_00000;
    timing4[3][4] = 16'b11001_100100_00000;
    timing4[3][5] = 16'b11111_111110_11111;
    timing4[3][6] = 16'b11111_111110_11111;
    timing4[3][7] = 16'b11111_111110_11111;
    timing4[3][8] = 16'b11111_111110_11111;
    timing4[3][9] = 16'b11111_111110_11111;
    timing4[3][10] = 16'b11001_100100_00000;
    timing4[3][11] = 16'b11111_101110_00000;
    timing4[3][12] = 16'b11111_101110_00000;
    timing4[3][13] = 16'b00000_000000_00000;
    timing4[3][14] = 16'b11111_111110_11111;
    timing4[4][0] = 16'b11111_111110_11111;
    timing4[4][1] = 16'b00000_000000_00000;
    timing4[4][2] = 16'b11111_101110_00000;
    timing4[4][3] = 16'b11001_100100_00000;
    timing4[4][4] = 16'b11111_111110_11111;
    timing4[4][5] = 16'b11111_111110_11111;
    timing4[4][6] = 16'b11111_111110_11111;
    timing4[4][7] = 16'b11111_111110_11111;
    timing4[4][8] = 16'b11111_111110_11111;
    timing4[4][9] = 16'b11111_111110_11111;
    timing4[4][10] = 16'b11111_111110_11111;
    timing4[4][11] = 16'b11001_100100_00000;
    timing4[4][12] = 16'b11111_101110_00000;
    timing4[4][13] = 16'b00000_000000_00000;
    timing4[4][14] = 16'b11111_111110_11111;
    timing4[5][0] = 16'b11111_111110_11111;
    timing4[5][1] = 16'b11111_101110_00000;
    timing4[5][2] = 16'b11001_100100_00000;
    timing4[5][3] = 16'b11111_111110_11111;
    timing4[5][4] = 16'b11111_111110_11111;
    timing4[5][5] = 16'b11111_111110_11111;
    timing4[5][6] = 16'b11111_111110_11111;
    timing4[5][7] = 16'b11111_111110_11111;
    timing4[5][8] = 16'b11111_111110_11111;
    timing4[5][9] = 16'b11111_111110_11111;
    timing4[5][10] = 16'b11111_111110_11111;
    timing4[5][11] = 16'b11111_111110_11111;
    timing4[5][12] = 16'b11001_100100_00000;
    timing4[5][13] = 16'b11111_101110_00000;
    timing4[5][14] = 16'b11111_111110_11111;
    timing4[6][0] = 16'b11111_111110_11111;
    timing4[6][1] = 16'b11111_101110_00000;
    timing4[6][2] = 16'b11001_100100_00000;
    timing4[6][3] = 16'b11111_111110_11111;
    timing4[6][4] = 16'b11111_111110_11111;
    timing4[6][5] = 16'b11111_111110_11111;
    timing4[6][6] = 16'b11111_111110_11111;
    timing4[6][7] = 16'b11111_111110_11111;
    timing4[6][8] = 16'b11111_111110_11111;
    timing4[6][9] = 16'b11111_111110_11111;
    timing4[6][10] = 16'b11111_111110_11111;
    timing4[6][11] = 16'b11111_111110_11111;
    timing4[6][12] = 16'b11001_100100_00000;
    timing4[6][13] = 16'b11111_101110_00000;
    timing4[6][14] = 16'b11111_111110_11111;
    timing4[7][0] = 16'b11111_111110_11111;
    timing4[7][1] = 16'b11111_101110_00000;
    timing4[7][2] = 16'b11001_100100_00000;
    timing4[7][3] = 16'b11111_111110_11111;
    timing4[7][4] = 16'b11111_111110_11111;
    timing4[7][5] = 16'b11111_111110_11111;
    timing4[7][6] = 16'b11111_111110_11111;
    timing4[7][7] = 16'b00000_000000_00000;
    timing4[7][8] = 16'b00000_000000_00000;
    timing4[7][9] = 16'b00000_000000_00000;
    timing4[7][10] = 16'b00000_000000_00000;
    timing4[7][11] = 16'b11111_111110_11111;
    timing4[7][12] = 16'b11001_100100_00000;
    timing4[7][13] = 16'b11111_101110_00000;
    timing4[7][14] = 16'b11111_111110_11111;
    timing4[8][0] = 16'b11111_111110_11111;
    timing4[8][1] = 16'b11111_101110_00000;
    timing4[8][2] = 16'b11001_100100_00000;
    timing4[8][3] = 16'b11111_111110_11111;
    timing4[8][4] = 16'b11111_111110_11111;
    timing4[8][5] = 16'b11111_111110_11111;
    timing4[8][6] = 16'b11111_111110_11111;
    timing4[8][7] = 16'b11111_111110_11111;
    timing4[8][8] = 16'b00111_001111_00111;
    timing4[8][9] = 16'b11111_111110_11111;
    timing4[8][10] = 16'b11111_111110_11111;
    timing4[8][11] = 16'b11111_111110_11111;
    timing4[8][12] = 16'b11001_100100_00000;
    timing4[8][13] = 16'b11111_101110_00000;
    timing4[8][14] = 16'b11111_111110_11111;
    timing4[9][0] = 16'b11111_111110_11111;
    timing4[9][1] = 16'b11111_101110_00000;
    timing4[9][2] = 16'b11001_100100_00000;
    timing4[9][3] = 16'b11111_111110_11111;
    timing4[9][4] = 16'b11111_111110_11111;
    timing4[9][5] = 16'b11111_111110_11111;
    timing4[9][6] = 16'b11111_111110_11111;
    timing4[9][7] = 16'b11111_111110_11111;
    timing4[9][8] = 16'b00111_001111_00111;
    timing4[9][9] = 16'b11111_111110_11111;
    timing4[9][10] = 16'b11111_111110_11111;
    timing4[9][11] = 16'b11111_111110_11111;
    timing4[9][12] = 16'b11001_100100_00000;
    timing4[9][13] = 16'b11111_101110_00000;
    timing4[9][14] = 16'b11111_111110_11111;
    timing4[10][0] = 16'b11111_111110_11111;
    timing4[10][1] = 16'b00000_000000_00000;
    timing4[10][2] = 16'b11111_101110_00000;
    timing4[10][3] = 16'b11001_100100_00000;
    timing4[10][4] = 16'b11111_111110_11111;
    timing4[10][5] = 16'b11111_111110_11111;
    timing4[10][6] = 16'b11111_111110_11111;
    timing4[10][7] = 16'b11111_111110_11111;
    timing4[10][8] = 16'b11111_111110_11111;
    timing4[10][9] = 16'b00111_001111_00111;
    timing4[10][10] = 16'b11111_111110_11111;
    timing4[10][11] = 16'b11001_100100_00000;
    timing4[10][12] = 16'b11111_101110_00000;
    timing4[10][13] = 16'b00000_000000_00000;
    timing4[10][14] = 16'b11111_111110_11111;
    timing4[11][0] = 16'b11111_111110_11111;
    timing4[11][1] = 16'b00000_000000_00000;
    timing4[11][2] = 16'b11111_101110_00000;
    timing4[11][3] = 16'b11111_101110_00000;
    timing4[11][4] = 16'b11001_100100_00000;
    timing4[11][5] = 16'b11111_111110_11111;
    timing4[11][6] = 16'b11111_111110_11111;
    timing4[11][7] = 16'b11111_111110_11111;
    timing4[11][8] = 16'b11111_111110_11111;
    timing4[11][9] = 16'b11111_111110_11111;
    timing4[11][10] = 16'b11001_100100_00000;
    timing4[11][11] = 16'b11111_101110_00000;
    timing4[11][12] = 16'b11111_101110_00000;
    timing4[11][13] = 16'b00000_000000_00000;
    timing4[11][14] = 16'b11111_111110_11111;
    timing4[12][0] = 16'b11111_111110_11111;
    timing4[12][1] = 16'b00000_000000_00000;
    timing4[12][2] = 16'b00000_000000_00000;
    timing4[12][3] = 16'b11111_101110_00000;
    timing4[12][4] = 16'b11111_101110_00000;
    timing4[12][5] = 16'b11001_100100_00000;
    timing4[12][6] = 16'b11001_100100_00000;
    timing4[12][7] = 16'b11001_100100_00000;
    timing4[12][8] = 16'b11001_100100_00000;
    timing4[12][9] = 16'b11001_100100_00000;
    timing4[12][10] = 16'b11111_101110_00000;
    timing4[12][11] = 16'b11111_101110_00000;
    timing4[12][12] = 16'b00000_000000_00000;
    timing4[12][13] = 16'b00000_000000_00000;
    timing4[12][14] = 16'b11111_111110_11111;
    timing4[13][0] = 16'b11111_111110_11111;
    timing4[13][1] = 16'b00000_000000_00000;
    timing4[13][2] = 16'b00000_000000_00000;
    timing4[13][3] = 16'b00000_000000_00000;
    timing4[13][4] = 16'b00000_000000_00000;
    timing4[13][5] = 16'b11111_101110_00000;
    timing4[13][6] = 16'b11111_101110_00000;
    timing4[13][7] = 16'b11111_101110_00000;
    timing4[13][8] = 16'b11111_101110_00000;
    timing4[13][9] = 16'b11111_101110_00000;
    timing4[13][10] = 16'b00000_000000_00000;
    timing4[13][11] = 16'b00000_000000_00000;
    timing4[13][12] = 16'b00000_000000_00000;
    timing4[13][13] = 16'b00000_000000_00000;
    timing4[13][14] = 16'b11111_111110_11111;
    timing4[14][0] = 16'b11111_111110_11111;
    timing4[14][1] = 16'b11111_111110_11111;
    timing4[14][2] = 16'b11111_111110_11111;
    timing4[14][3] = 16'b11111_111110_11111;
    timing4[14][4] = 16'b11111_111110_11111;
    timing4[14][5] = 16'b11111_111110_11111;
    timing4[14][6] = 16'b11111_111110_11111;
    timing4[14][7] = 16'b11111_111110_11111;
    timing4[14][8] = 16'b11111_111110_11111;
    timing4[14][9] = 16'b11111_111110_11111;
    timing4[14][10] = 16'b11111_111110_11111;
    timing4[14][11] = 16'b11111_111110_11111;
    timing4[14][12] = 16'b11111_111110_11111;
    timing4[14][13] = 16'b11111_111110_11111;
    timing4[14][14] = 16'b11111_111110_11111;
    
    timing5[0][0] = 16'b11111_111110_11111;
    timing5[0][1] = 16'b11111_111110_11111;
    timing5[0][2] = 16'b11111_111110_11111;
    timing5[0][3] = 16'b11111_111110_11111;
    timing5[0][4] = 16'b11111_111110_11111;
    timing5[0][5] = 16'b11111_111110_11111;
    timing5[0][6] = 16'b11111_111110_11111;
    timing5[0][7] = 16'b11111_111110_11111;
    timing5[0][8] = 16'b11111_111110_11111;
    timing5[0][9] = 16'b11111_111110_11111;
    timing5[0][10] = 16'b11111_111110_11111;
    timing5[0][11] = 16'b11111_111110_11111;
    timing5[0][12] = 16'b11111_111110_11111;
    timing5[0][13] = 16'b11111_111110_11111;
    timing5[0][14] = 16'b11111_111110_11111;
    timing5[1][0] = 16'b11111_111110_11111;
    timing5[1][1] = 16'b00000_000000_00000;
    timing5[1][2] = 16'b00000_000000_00000;
    timing5[1][3] = 16'b00000_000000_00000;
    timing5[1][4] = 16'b00000_000000_00000;
    timing5[1][5] = 16'b11111_101110_00000;
    timing5[1][6] = 16'b11111_101110_00000;
    timing5[1][7] = 16'b11111_101110_00000;
    timing5[1][8] = 16'b11111_101110_00000;
    timing5[1][9] = 16'b11111_101110_00000;
    timing5[1][10] = 16'b00000_000000_00000;
    timing5[1][11] = 16'b00000_000000_00000;
    timing5[1][12] = 16'b00000_000000_00000;
    timing5[1][13] = 16'b00000_000000_00000;
    timing5[1][14] = 16'b11111_111110_11111;
    timing5[2][0] = 16'b11111_111110_11111;
    timing5[2][1] = 16'b00000_000000_00000;
    timing5[2][2] = 16'b00000_000000_00000;
    timing5[2][3] = 16'b11111_101110_00000;
    timing5[2][4] = 16'b11111_101110_00000;
    timing5[2][5] = 16'b11001_100100_00000;
    timing5[2][6] = 16'b11001_100100_00000;
    timing5[2][7] = 16'b11001_100100_00000;
    timing5[2][8] = 16'b11001_100100_00000;
    timing5[2][9] = 16'b11001_100100_00000;
    timing5[2][10] = 16'b11111_101110_00000;
    timing5[2][11] = 16'b11111_101110_00000;
    timing5[2][12] = 16'b00000_000000_00000;
    timing5[2][13] = 16'b00000_000000_00000;
    timing5[2][14] = 16'b11111_111110_11111;
    timing5[3][0] = 16'b11111_111110_11111;
    timing5[3][1] = 16'b00000_000000_00000;
    timing5[3][2] = 16'b11111_101110_00000;
    timing5[3][3] = 16'b11111_101110_00000;
    timing5[3][4] = 16'b11001_100100_00000;
    timing5[3][5] = 16'b11111_111110_11111;
    timing5[3][6] = 16'b11111_111110_11111;
    timing5[3][7] = 16'b11111_111110_11111;
    timing5[3][8] = 16'b11111_111110_11111;
    timing5[3][9] = 16'b11111_111110_11111;
    timing5[3][10] = 16'b11001_100100_00000;
    timing5[3][11] = 16'b11111_101110_00000;
    timing5[3][12] = 16'b11111_101110_00000;
    timing5[3][13] = 16'b00000_000000_00000;
    timing5[3][14] = 16'b11111_111110_11111;
    timing5[4][0] = 16'b11111_111110_11111;
    timing5[4][1] = 16'b00000_000000_00000;
    timing5[4][2] = 16'b11111_101110_00000;
    timing5[4][3] = 16'b11001_100100_00000;
    timing5[4][4] = 16'b11111_111110_11111;
    timing5[4][5] = 16'b11111_111110_11111;
    timing5[4][6] = 16'b11111_111110_11111;
    timing5[4][7] = 16'b11111_111110_11111;
    timing5[4][8] = 16'b11111_111110_11111;
    timing5[4][9] = 16'b11111_111110_11111;
    timing5[4][10] = 16'b11111_111110_11111;
    timing5[4][11] = 16'b11001_100100_00000;
    timing5[4][12] = 16'b11111_101110_00000;
    timing5[4][13] = 16'b00000_000000_00000;
    timing5[4][14] = 16'b11111_111110_11111;
    timing5[5][0] = 16'b11111_111110_11111;
    timing5[5][1] = 16'b11111_101110_00000;
    timing5[5][2] = 16'b11001_100100_00000;
    timing5[5][3] = 16'b11111_111110_11111;
    timing5[5][4] = 16'b11111_111110_11111;
    timing5[5][5] = 16'b11111_111110_11111;
    timing5[5][6] = 16'b11111_111110_11111;
    timing5[5][7] = 16'b11111_111110_11111;
    timing5[5][8] = 16'b11111_111110_11111;
    timing5[5][9] = 16'b11111_111110_11111;
    timing5[5][10] = 16'b11111_111110_11111;
    timing5[5][11] = 16'b11111_111110_11111;
    timing5[5][12] = 16'b11001_100100_00000;
    timing5[5][13] = 16'b11111_101110_00000;
    timing5[5][14] = 16'b11111_111110_11111;
    timing5[6][0] = 16'b11111_111110_11111;
    timing5[6][1] = 16'b11111_101110_00000;
    timing5[6][2] = 16'b11001_100100_00000;
    timing5[6][3] = 16'b11111_111110_11111;
    timing5[6][4] = 16'b11111_111110_11111;
    timing5[6][5] = 16'b11111_111110_11111;
    timing5[6][6] = 16'b11111_111110_11111;
    timing5[6][7] = 16'b11111_111110_11111;
    timing5[6][8] = 16'b11111_111110_11111;
    timing5[6][9] = 16'b11111_111110_11111;
    timing5[6][10] = 16'b11111_111110_11111;
    timing5[6][11] = 16'b11111_111110_11111;
    timing5[6][12] = 16'b11001_100100_00000;
    timing5[6][13] = 16'b11111_101110_00000;
    timing5[6][14] = 16'b11111_111110_11111;
    timing5[7][0] = 16'b11111_111110_11111;
    timing5[7][1] = 16'b11111_101110_00000;
    timing5[7][2] = 16'b11001_100100_00000;
    timing5[7][3] = 16'b11111_111110_11111;
    timing5[7][4] = 16'b11111_111110_11111;
    timing5[7][5] = 16'b11111_111110_11111;
    timing5[7][6] = 16'b11111_111110_11111;
    timing5[7][7] = 16'b00000_000000_00000;
    timing5[7][8] = 16'b00000_000000_00000;
    timing5[7][9] = 16'b00000_000000_00000;
    timing5[7][10] = 16'b00000_000000_00000;
    timing5[7][11] = 16'b11111_111110_11111;
    timing5[7][12] = 16'b11001_100100_00000;
    timing5[7][13] = 16'b11111_101110_00000;
    timing5[7][14] = 16'b11111_111110_11111;
    timing5[8][0] = 16'b11111_111110_11111;
    timing5[8][1] = 16'b11111_101110_00000;
    timing5[8][2] = 16'b11001_100100_00000;
    timing5[8][3] = 16'b11111_111110_11111;
    timing5[8][4] = 16'b11111_111110_11111;
    timing5[8][5] = 16'b11111_111110_11111;
    timing5[8][6] = 16'b11111_111110_11111;
    timing5[8][7] = 16'b00111_001111_00111;
    timing5[8][8] = 16'b11111_111110_11111;
    timing5[8][9] = 16'b11111_111110_11111;
    timing5[8][10] = 16'b11111_111110_11111;
    timing5[8][11] = 16'b11111_111110_11111;
    timing5[8][12] = 16'b11001_100100_00000;
    timing5[8][13] = 16'b11111_101110_00000;
    timing5[8][14] = 16'b11111_111110_11111;
    timing5[9][0] = 16'b11111_111110_11111;
    timing5[9][1] = 16'b11111_101110_00000;
    timing5[9][2] = 16'b11001_100100_00000;
    timing5[9][3] = 16'b11111_111110_11111;
    timing5[9][4] = 16'b11111_111110_11111;
    timing5[9][5] = 16'b11111_111110_11111;
    timing5[9][6] = 16'b11111_111110_11111;
    timing5[9][7] = 16'b00111_001111_00111;
    timing5[9][8] = 16'b11111_111110_11111;
    timing5[9][9] = 16'b11111_111110_11111;
    timing5[9][10] = 16'b11111_111110_11111;
    timing5[9][11] = 16'b11111_111110_11111;
    timing5[9][12] = 16'b11001_100100_00000;
    timing5[9][13] = 16'b11111_101110_00000;
    timing5[9][14] = 16'b11111_111110_11111;
    timing5[10][0] = 16'b11111_111110_11111;
    timing5[10][1] = 16'b00000_000000_00000;
    timing5[10][2] = 16'b11111_101110_00000;
    timing5[10][3] = 16'b11001_100100_00000;
    timing5[10][4] = 16'b11111_111110_11111;
    timing5[10][5] = 16'b11111_111110_11111;
    timing5[10][6] = 16'b11111_111110_11111;
    timing5[10][7] = 16'b00111_001111_00111;
    timing5[10][8] = 16'b11111_111110_11111;
    timing5[10][9] = 16'b11111_111110_11111;
    timing5[10][10] = 16'b11111_111110_11111;
    timing5[10][11] = 16'b11001_100100_00000;
    timing5[10][12] = 16'b11111_101110_00000;
    timing5[10][13] = 16'b00000_000000_00000;
    timing5[10][14] = 16'b11111_111110_11111;
    timing5[11][0] = 16'b11111_111110_11111;
    timing5[11][1] = 16'b00000_000000_00000;
    timing5[11][2] = 16'b11111_101110_00000;
    timing5[11][3] = 16'b11111_101110_00000;
    timing5[11][4] = 16'b11001_100100_00000;
    timing5[11][5] = 16'b11111_111110_11111;
    timing5[11][6] = 16'b11111_111110_11111;
    timing5[11][7] = 16'b00111_001111_00111;
    timing5[11][8] = 16'b11111_111110_11111;
    timing5[11][9] = 16'b11111_111110_11111;
    timing5[11][10] = 16'b11001_100100_00000;
    timing5[11][11] = 16'b11111_101110_00000;
    timing5[11][12] = 16'b11111_101110_00000;
    timing5[11][13] = 16'b00000_000000_00000;
    timing5[11][14] = 16'b11111_111110_11111;
    timing5[12][0] = 16'b11111_111110_11111;
    timing5[12][1] = 16'b00000_000000_00000;
    timing5[12][2] = 16'b00000_000000_00000;
    timing5[12][3] = 16'b11111_101110_00000;
    timing5[12][4] = 16'b11111_101110_00000;
    timing5[12][5] = 16'b11001_100100_00000;
    timing5[12][6] = 16'b11001_100100_00000;
    timing5[12][7] = 16'b11001_100100_00000;
    timing5[12][8] = 16'b11001_100100_00000;
    timing5[12][9] = 16'b11001_100100_00000;
    timing5[12][10] = 16'b11111_101110_00000;
    timing5[12][11] = 16'b11111_101110_00000;
    timing5[12][12] = 16'b00000_000000_00000;
    timing5[12][13] = 16'b00000_000000_00000;
    timing5[12][14] = 16'b11111_111110_11111;
    timing5[13][0] = 16'b11111_111110_11111;
    timing5[13][1] = 16'b00000_000000_00000;
    timing5[13][2] = 16'b00000_000000_00000;
    timing5[13][3] = 16'b00000_000000_00000;
    timing5[13][4] = 16'b00000_000000_00000;
    timing5[13][5] = 16'b11111_101110_00000;
    timing5[13][6] = 16'b11111_101110_00000;
    timing5[13][7] = 16'b11111_101110_00000;
    timing5[13][8] = 16'b11111_101110_00000;
    timing5[13][9] = 16'b11111_101110_00000;
    timing5[13][10] = 16'b00000_000000_00000;
    timing5[13][11] = 16'b00000_000000_00000;
    timing5[13][12] = 16'b00000_000000_00000;
    timing5[13][13] = 16'b00000_000000_00000;
    timing5[13][14] = 16'b11111_111110_11111;
    timing5[14][0] = 16'b11111_111110_11111;
    timing5[14][1] = 16'b11111_111110_11111;
    timing5[14][2] = 16'b11111_111110_11111;
    timing5[14][3] = 16'b11111_111110_11111;
    timing5[14][4] = 16'b11111_111110_11111;
    timing5[14][5] = 16'b11111_111110_11111;
    timing5[14][6] = 16'b11111_111110_11111;
    timing5[14][7] = 16'b11111_111110_11111;
    timing5[14][8] = 16'b11111_111110_11111;
    timing5[14][9] = 16'b11111_111110_11111;
    timing5[14][10] = 16'b11111_111110_11111;
    timing5[14][11] = 16'b11111_111110_11111;
    timing5[14][12] = 16'b11111_111110_11111;
    timing5[14][13] = 16'b11111_111110_11111;
    timing5[14][14] = 16'b11111_111110_11111;
    
    timing6[0][0] = 16'b11111_111110_11111;
    timing6[0][1] = 16'b11111_111110_11111;
    timing6[0][2] = 16'b11111_111110_11111;
    timing6[0][3] = 16'b11111_111110_11111;
    timing6[0][4] = 16'b11111_111110_11111;
    timing6[0][5] = 16'b11111_111110_11111;
    timing6[0][6] = 16'b11111_111110_11111;
    timing6[0][7] = 16'b11111_111110_11111;
    timing6[0][8] = 16'b11111_111110_11111;
    timing6[0][9] = 16'b11111_111110_11111;
    timing6[0][10] = 16'b11111_111110_11111;
    timing6[0][11] = 16'b11111_111110_11111;
    timing6[0][12] = 16'b11111_111110_11111;
    timing6[0][13] = 16'b11111_111110_11111;
    timing6[0][14] = 16'b11111_111110_11111;
    timing6[1][0] = 16'b11111_111110_11111;
    timing6[1][1] = 16'b00000_000000_00000;
    timing6[1][2] = 16'b00000_000000_00000;
    timing6[1][3] = 16'b00000_000000_00000;
    timing6[1][4] = 16'b00000_000000_00000;
    timing6[1][5] = 16'b11111_101110_00000;
    timing6[1][6] = 16'b11111_101110_00000;
    timing6[1][7] = 16'b11111_101110_00000;
    timing6[1][8] = 16'b11111_101110_00000;
    timing6[1][9] = 16'b11111_101110_00000;
    timing6[1][10] = 16'b00000_000000_00000;
    timing6[1][11] = 16'b00000_000000_00000;
    timing6[1][12] = 16'b00000_000000_00000;
    timing6[1][13] = 16'b00000_000000_00000;
    timing6[1][14] = 16'b11111_111110_11111;
    timing6[2][0] = 16'b11111_111110_11111;
    timing6[2][1] = 16'b00000_000000_00000;
    timing6[2][2] = 16'b00000_000000_00000;
    timing6[2][3] = 16'b11111_101110_00000;
    timing6[2][4] = 16'b11111_101110_00000;
    timing6[2][5] = 16'b11001_100100_00000;
    timing6[2][6] = 16'b11001_100100_00000;
    timing6[2][7] = 16'b11001_100100_00000;
    timing6[2][8] = 16'b11001_100100_00000;
    timing6[2][9] = 16'b11001_100100_00000;
    timing6[2][10] = 16'b11111_101110_00000;
    timing6[2][11] = 16'b11111_101110_00000;
    timing6[2][12] = 16'b00000_000000_00000;
    timing6[2][13] = 16'b00000_000000_00000;
    timing6[2][14] = 16'b11111_111110_11111;
    timing6[3][0] = 16'b11111_111110_11111;
    timing6[3][1] = 16'b00000_000000_00000;
    timing6[3][2] = 16'b11111_101110_00000;
    timing6[3][3] = 16'b11111_101110_00000;
    timing6[3][4] = 16'b11001_100100_00000;
    timing6[3][5] = 16'b11111_111110_11111;
    timing6[3][6] = 16'b11111_111110_11111;
    timing6[3][7] = 16'b11111_111110_11111;
    timing6[3][8] = 16'b11111_111110_11111;
    timing6[3][9] = 16'b11111_111110_11111;
    timing6[3][10] = 16'b11001_100100_00000;
    timing6[3][11] = 16'b11111_101110_00000;
    timing6[3][12] = 16'b11111_101110_00000;
    timing6[3][13] = 16'b00000_000000_00000;
    timing6[3][14] = 16'b11111_111110_11111;
    timing6[4][0] = 16'b11111_111110_11111;
    timing6[4][1] = 16'b00000_000000_00000;
    timing6[4][2] = 16'b11111_101110_00000;
    timing6[4][3] = 16'b11001_100100_00000;
    timing6[4][4] = 16'b11111_111110_11111;
    timing6[4][5] = 16'b11111_111110_11111;
    timing6[4][6] = 16'b11111_111110_11111;
    timing6[4][7] = 16'b11111_111110_11111;
    timing6[4][8] = 16'b11111_111110_11111;
    timing6[4][9] = 16'b11111_111110_11111;
    timing6[4][10] = 16'b11111_111110_11111;
    timing6[4][11] = 16'b11001_100100_00000;
    timing6[4][12] = 16'b11111_101110_00000;
    timing6[4][13] = 16'b00000_000000_00000;
    timing6[4][14] = 16'b11111_111110_11111;
    timing6[5][0] = 16'b11111_111110_11111;
    timing6[5][1] = 16'b11111_101110_00000;
    timing6[5][2] = 16'b11001_100100_00000;
    timing6[5][3] = 16'b11111_111110_11111;
    timing6[5][4] = 16'b11111_111110_11111;
    timing6[5][5] = 16'b11111_111110_11111;
    timing6[5][6] = 16'b11111_111110_11111;
    timing6[5][7] = 16'b11111_111110_11111;
    timing6[5][8] = 16'b11111_111110_11111;
    timing6[5][9] = 16'b11111_111110_11111;
    timing6[5][10] = 16'b11111_111110_11111;
    timing6[5][11] = 16'b11111_111110_11111;
    timing6[5][12] = 16'b11001_100100_00000;
    timing6[5][13] = 16'b11111_101110_00000;
    timing6[5][14] = 16'b11111_111110_11111;
    timing6[6][0] = 16'b11111_111110_11111;
    timing6[6][1] = 16'b11111_101110_00000;
    timing6[6][2] = 16'b11001_100100_00000;
    timing6[6][3] = 16'b11111_111110_11111;
    timing6[6][4] = 16'b11111_111110_11111;
    timing6[6][5] = 16'b11111_111110_11111;
    timing6[6][6] = 16'b11111_111110_11111;
    timing6[6][7] = 16'b11111_111110_11111;
    timing6[6][8] = 16'b11111_111110_11111;
    timing6[6][9] = 16'b11111_111110_11111;
    timing6[6][10] = 16'b11111_111110_11111;
    timing6[6][11] = 16'b11111_111110_11111;
    timing6[6][12] = 16'b11001_100100_00000;
    timing6[6][13] = 16'b11111_101110_00000;
    timing6[6][14] = 16'b11111_111110_11111;
    timing6[7][0] = 16'b11111_111110_11111;
    timing6[7][1] = 16'b11111_101110_00000;
    timing6[7][2] = 16'b11001_100100_00000;
    timing6[7][3] = 16'b11111_111110_11111;
    timing6[7][4] = 16'b11111_111110_11111;
    timing6[7][5] = 16'b11111_111110_11111;
    timing6[7][6] = 16'b11111_111110_11111;
    timing6[7][7] = 16'b00000_000000_00000;
    timing6[7][8] = 16'b00000_000000_00000;
    timing6[7][9] = 16'b00000_000000_00000;
    timing6[7][10] = 16'b00000_000000_00000;
    timing6[7][11] = 16'b11111_111110_11111;
    timing6[7][12] = 16'b11001_100100_00000;
    timing6[7][13] = 16'b11111_101110_00000;
    timing6[7][14] = 16'b11111_111110_11111;
    timing6[8][0] = 16'b11111_111110_11111;
    timing6[8][1] = 16'b11111_101110_00000;
    timing6[8][2] = 16'b11001_100100_00000;
    timing6[8][3] = 16'b11111_111110_11111;
    timing6[8][4] = 16'b11111_111110_11111;
    timing6[8][5] = 16'b11111_111110_11111;
    timing6[8][6] = 16'b00111_001111_00111;
    timing6[8][7] = 16'b11111_111110_11111;
    timing6[8][8] = 16'b11111_111110_11111;
    timing6[8][9] = 16'b11111_111110_11111;
    timing6[8][10] = 16'b11111_111110_11111;
    timing6[8][11] = 16'b11111_111110_11111;
    timing6[8][12] = 16'b11001_100100_00000;
    timing6[8][13] = 16'b11111_101110_00000;
    timing6[8][14] = 16'b11111_111110_11111;
    timing6[9][0] = 16'b11111_111110_11111;
    timing6[9][1] = 16'b11111_101110_00000;
    timing6[9][2] = 16'b11001_100100_00000;
    timing6[9][3] = 16'b11111_111110_11111;
    timing6[9][4] = 16'b11111_111110_11111;
    timing6[9][5] = 16'b00111_001111_00111;
    timing6[9][6] = 16'b11111_111110_11111;
    timing6[9][7] = 16'b11111_111110_11111;
    timing6[9][8] = 16'b11111_111110_11111;
    timing6[9][9] = 16'b11111_111110_11111;
    timing6[9][10] = 16'b11111_111110_11111;
    timing6[9][11] = 16'b11111_111110_11111;
    timing6[9][12] = 16'b11001_100100_00000;
    timing6[9][13] = 16'b11111_101110_00000;
    timing6[9][14] = 16'b11111_111110_11111;
    timing6[10][0] = 16'b11111_111110_11111;
    timing6[10][1] = 16'b00000_000000_00000;
    timing6[10][2] = 16'b11111_101110_00000;
    timing6[10][3] = 16'b11001_100100_00000;
    timing6[10][4] = 16'b11111_111110_11111;
    timing6[10][5] = 16'b00111_001111_00111;
    timing6[10][6] = 16'b11111_111110_11111;
    timing6[10][7] = 16'b11111_111110_11111;
    timing6[10][8] = 16'b11111_111110_11111;
    timing6[10][9] = 16'b11111_111110_11111;
    timing6[10][10] = 16'b11111_111110_11111;
    timing6[10][11] = 16'b11001_100100_00000;
    timing6[10][12] = 16'b11111_101110_00000;
    timing6[10][13] = 16'b00000_000000_00000;
    timing6[10][14] = 16'b11111_111110_11111;
    timing6[11][0] = 16'b11111_111110_11111;
    timing6[11][1] = 16'b00000_000000_00000;
    timing6[11][2] = 16'b11111_101110_00000;
    timing6[11][3] = 16'b11111_101110_00000;
    timing6[11][4] = 16'b11001_100100_00000;
    timing6[11][5] = 16'b11111_111110_11111;
    timing6[11][6] = 16'b11111_111110_11111;
    timing6[11][7] = 16'b11111_111110_11111;
    timing6[11][8] = 16'b11111_111110_11111;
    timing6[11][9] = 16'b11111_111110_11111;
    timing6[11][10] = 16'b11001_100100_00000;
    timing6[11][11] = 16'b11111_101110_00000;
    timing6[11][12] = 16'b11111_101110_00000;
    timing6[11][13] = 16'b00000_000000_00000;
    timing6[11][14] = 16'b11111_111110_11111;
    timing6[12][0] = 16'b11111_111110_11111;
    timing6[12][1] = 16'b00000_000000_00000;
    timing6[12][2] = 16'b00000_000000_00000;
    timing6[12][3] = 16'b11111_101110_00000;
    timing6[12][4] = 16'b11111_101110_00000;
    timing6[12][5] = 16'b11001_100100_00000;
    timing6[12][6] = 16'b11001_100100_00000;
    timing6[12][7] = 16'b11001_100100_00000;
    timing6[12][8] = 16'b11001_100100_00000;
    timing6[12][9] = 16'b11001_100100_00000;
    timing6[12][10] = 16'b11111_101110_00000;
    timing6[12][11] = 16'b11111_101110_00000;
    timing6[12][12] = 16'b00000_000000_00000;
    timing6[12][13] = 16'b00000_000000_00000;
    timing6[12][14] = 16'b11111_111110_11111;
    timing6[13][0] = 16'b11111_111110_11111;
    timing6[13][1] = 16'b00000_000000_00000;
    timing6[13][2] = 16'b00000_000000_00000;
    timing6[13][3] = 16'b00000_000000_00000;
    timing6[13][4] = 16'b00000_000000_00000;
    timing6[13][5] = 16'b11111_101110_00000;
    timing6[13][6] = 16'b11111_101110_00000;
    timing6[13][7] = 16'b11111_101110_00000;
    timing6[13][8] = 16'b11111_101110_00000;
    timing6[13][9] = 16'b11111_101110_00000;
    timing6[13][10] = 16'b00000_000000_00000;
    timing6[13][11] = 16'b00000_000000_00000;
    timing6[13][12] = 16'b00000_000000_00000;
    timing6[13][13] = 16'b00000_000000_00000;
    timing6[13][14] = 16'b11111_111110_11111;
    timing6[14][0] = 16'b11111_111110_11111;
    timing6[14][1] = 16'b11111_111110_11111;
    timing6[14][2] = 16'b11111_111110_11111;
    timing6[14][3] = 16'b11111_111110_11111;
    timing6[14][4] = 16'b11111_111110_11111;
    timing6[14][5] = 16'b11111_111110_11111;
    timing6[14][6] = 16'b11111_111110_11111;
    timing6[14][7] = 16'b11111_111110_11111;
    timing6[14][8] = 16'b11111_111110_11111;
    timing6[14][9] = 16'b11111_111110_11111;
    timing6[14][10] = 16'b11111_111110_11111;
    timing6[14][11] = 16'b11111_111110_11111;
    timing6[14][12] = 16'b11111_111110_11111;
    timing6[14][13] = 16'b11111_111110_11111;
    timing6[14][14] = 16'b11111_111110_11111;
    
    timing7[0][0] = 16'b11111_111110_11111;
    timing7[0][1] = 16'b11111_111110_11111;
    timing7[0][2] = 16'b11111_111110_11111;
    timing7[0][3] = 16'b11111_111110_11111;
    timing7[0][4] = 16'b11111_111110_11111;
    timing7[0][5] = 16'b11111_111110_11111;
    timing7[0][6] = 16'b11111_111110_11111;
    timing7[0][7] = 16'b11111_111110_11111;
    timing7[0][8] = 16'b11111_111110_11111;
    timing7[0][9] = 16'b11111_111110_11111;
    timing7[0][10] = 16'b11111_111110_11111;
    timing7[0][11] = 16'b11111_111110_11111;
    timing7[0][12] = 16'b11111_111110_11111;
    timing7[0][13] = 16'b11111_111110_11111;
    timing7[0][14] = 16'b11111_111110_11111;
    timing7[1][0] = 16'b11111_111110_11111;
    timing7[1][1] = 16'b00000_000000_00000;
    timing7[1][2] = 16'b00000_000000_00000;
    timing7[1][3] = 16'b00000_000000_00000;
    timing7[1][4] = 16'b00000_000000_00000;
    timing7[1][5] = 16'b11111_101110_00000;
    timing7[1][6] = 16'b11111_101110_00000;
    timing7[1][7] = 16'b11111_101110_00000;
    timing7[1][8] = 16'b11111_101110_00000;
    timing7[1][9] = 16'b11111_101110_00000;
    timing7[1][10] = 16'b00000_000000_00000;
    timing7[1][11] = 16'b00000_000000_00000;
    timing7[1][12] = 16'b00000_000000_00000;
    timing7[1][13] = 16'b00000_000000_00000;
    timing7[1][14] = 16'b11111_111110_11111;
    timing7[2][0] = 16'b11111_111110_11111;
    timing7[2][1] = 16'b00000_000000_00000;
    timing7[2][2] = 16'b00000_000000_00000;
    timing7[2][3] = 16'b11111_101110_00000;
    timing7[2][4] = 16'b11111_101110_00000;
    timing7[2][5] = 16'b11001_100100_00000;
    timing7[2][6] = 16'b11001_100100_00000;
    timing7[2][7] = 16'b11001_100100_00000;
    timing7[2][8] = 16'b11001_100100_00000;
    timing7[2][9] = 16'b11001_100100_00000;
    timing7[2][10] = 16'b11111_101110_00000;
    timing7[2][11] = 16'b11111_101110_00000;
    timing7[2][12] = 16'b00000_000000_00000;
    timing7[2][13] = 16'b00000_000000_00000;
    timing7[2][14] = 16'b11111_111110_11111;
    timing7[3][0] = 16'b11111_111110_11111;
    timing7[3][1] = 16'b00000_000000_00000;
    timing7[3][2] = 16'b11111_101110_00000;
    timing7[3][3] = 16'b11111_101110_00000;
    timing7[3][4] = 16'b11001_100100_00000;
    timing7[3][5] = 16'b11111_111110_11111;
    timing7[3][6] = 16'b11111_111110_11111;
    timing7[3][7] = 16'b11111_111110_11111;
    timing7[3][8] = 16'b11111_111110_11111;
    timing7[3][9] = 16'b11111_111110_11111;
    timing7[3][10] = 16'b11001_100100_00000;
    timing7[3][11] = 16'b11111_101110_00000;
    timing7[3][12] = 16'b11111_101110_00000;
    timing7[3][13] = 16'b00000_000000_00000;
    timing7[3][14] = 16'b11111_111110_11111;
    timing7[4][0] = 16'b11111_111110_11111;
    timing7[4][1] = 16'b00000_000000_00000;
    timing7[4][2] = 16'b11111_101110_00000;
    timing7[4][3] = 16'b11001_100100_00000;
    timing7[4][4] = 16'b11111_111110_11111;
    timing7[4][5] = 16'b11111_111110_11111;
    timing7[4][6] = 16'b11111_111110_11111;
    timing7[4][7] = 16'b11111_111110_11111;
    timing7[4][8] = 16'b11111_111110_11111;
    timing7[4][9] = 16'b11111_111110_11111;
    timing7[4][10] = 16'b11111_111110_11111;
    timing7[4][11] = 16'b11001_100100_00000;
    timing7[4][12] = 16'b11111_101110_00000;
    timing7[4][13] = 16'b00000_000000_00000;
    timing7[4][14] = 16'b11111_111110_11111;
    timing7[5][0] = 16'b11111_111110_11111;
    timing7[5][1] = 16'b11111_101110_00000;
    timing7[5][2] = 16'b11001_100100_00000;
    timing7[5][3] = 16'b11111_111110_11111;
    timing7[5][4] = 16'b11111_111110_11111;
    timing7[5][5] = 16'b11111_111110_11111;
    timing7[5][6] = 16'b11111_111110_11111;
    timing7[5][7] = 16'b11111_111110_11111;
    timing7[5][8] = 16'b11111_111110_11111;
    timing7[5][9] = 16'b11111_111110_11111;
    timing7[5][10] = 16'b11111_111110_11111;
    timing7[5][11] = 16'b11111_111110_11111;
    timing7[5][12] = 16'b11001_100100_00000;
    timing7[5][13] = 16'b11111_101110_00000;
    timing7[5][14] = 16'b11111_111110_11111;
    timing7[6][0] = 16'b11111_111110_11111;
    timing7[6][1] = 16'b11111_101110_00000;
    timing7[6][2] = 16'b11001_100100_00000;
    timing7[6][3] = 16'b11111_111110_11111;
    timing7[6][4] = 16'b11111_111110_11111;
    timing7[6][5] = 16'b11111_111110_11111;
    timing7[6][6] = 16'b11111_111110_11111;
    timing7[6][7] = 16'b11111_111110_11111;
    timing7[6][8] = 16'b11111_111110_11111;
    timing7[6][9] = 16'b11111_111110_11111;
    timing7[6][10] = 16'b11111_111110_11111;
    timing7[6][11] = 16'b11111_111110_11111;
    timing7[6][12] = 16'b11001_100100_00000;
    timing7[6][13] = 16'b11111_101110_00000;
    timing7[6][14] = 16'b11111_111110_11111;
    timing7[7][0] = 16'b11111_111110_11111;
    timing7[7][1] = 16'b11111_101110_00000;
    timing7[7][2] = 16'b11001_100100_00000;
    timing7[7][3] = 16'b00111_001111_00111;
    timing7[7][4] = 16'b00111_001111_00111;
    timing7[7][5] = 16'b00111_001111_00111;
    timing7[7][6] = 16'b00111_001111_00111;
    timing7[7][7] = 16'b00000_000000_00000;
    timing7[7][8] = 16'b00000_000000_00000;
    timing7[7][9] = 16'b00000_000000_00000;
    timing7[7][10] = 16'b00000_000000_00000;
    timing7[7][11] = 16'b11111_111110_11111;
    timing7[7][12] = 16'b11001_100100_00000;
    timing7[7][13] = 16'b11111_101110_00000;
    timing7[7][14] = 16'b11111_111110_11111;
    timing7[8][0] = 16'b11111_111110_11111;
    timing7[8][1] = 16'b11111_101110_00000;
    timing7[8][2] = 16'b11001_100100_00000;
    timing7[8][3] = 16'b11111_111110_11111;
    timing7[8][4] = 16'b11111_111110_11111;
    timing7[8][5] = 16'b11111_111110_11111;
    timing7[8][6] = 16'b11111_111110_11111;
    timing7[8][7] = 16'b11111_111110_11111;
    timing7[8][8] = 16'b11111_111110_11111;
    timing7[8][9] = 16'b11111_111110_11111;
    timing7[8][10] = 16'b11111_111110_11111;
    timing7[8][11] = 16'b11111_111110_11111;
    timing7[8][12] = 16'b11001_100100_00000;
    timing7[8][13] = 16'b11111_101110_00000;
    timing7[8][14] = 16'b11111_111110_11111;
    timing7[9][0] = 16'b11111_111110_11111;
    timing7[9][1] = 16'b11111_101110_00000;
    timing7[9][2] = 16'b11001_100100_00000;
    timing7[9][3] = 16'b11111_111110_11111;
    timing7[9][4] = 16'b11111_111110_11111;
    timing7[9][5] = 16'b11111_111110_11111;
    timing7[9][6] = 16'b11111_111110_11111;
    timing7[9][7] = 16'b11111_111110_11111;
    timing7[9][8] = 16'b11111_111110_11111;
    timing7[9][9] = 16'b11111_111110_11111;
    timing7[9][10] = 16'b11111_111110_11111;
    timing7[9][11] = 16'b11111_111110_11111;
    timing7[9][12] = 16'b11001_100100_00000;
    timing7[9][13] = 16'b11111_101110_00000;
    timing7[9][14] = 16'b11111_111110_11111;
    timing7[10][0] = 16'b11111_111110_11111;
    timing7[10][1] = 16'b00000_000000_00000;
    timing7[10][2] = 16'b11111_101110_00000;
    timing7[10][3] = 16'b11001_100100_00000;
    timing7[10][4] = 16'b11111_111110_11111;
    timing7[10][5] = 16'b11111_111110_11111;
    timing7[10][6] = 16'b11111_111110_11111;
    timing7[10][7] = 16'b11111_111110_11111;
    timing7[10][8] = 16'b11111_111110_11111;
    timing7[10][9] = 16'b11111_111110_11111;
    timing7[10][10] = 16'b11111_111110_11111;
    timing7[10][11] = 16'b11001_100100_00000;
    timing7[10][12] = 16'b11111_101110_00000;
    timing7[10][13] = 16'b00000_000000_00000;
    timing7[10][14] = 16'b11111_111110_11111;
    timing7[11][0] = 16'b11111_111110_11111;
    timing7[11][1] = 16'b00000_000000_00000;
    timing7[11][2] = 16'b11111_101110_00000;
    timing7[11][3] = 16'b11111_101110_00000;
    timing7[11][4] = 16'b11001_100100_00000;
    timing7[11][5] = 16'b11111_111110_11111;
    timing7[11][6] = 16'b11111_111110_11111;
    timing7[11][7] = 16'b11111_111110_11111;
    timing7[11][8] = 16'b11111_111110_11111;
    timing7[11][9] = 16'b11111_111110_11111;
    timing7[11][10] = 16'b11001_100100_00000;
    timing7[11][11] = 16'b11111_101110_00000;
    timing7[11][12] = 16'b11111_101110_00000;
    timing7[11][13] = 16'b00000_000000_00000;
    timing7[11][14] = 16'b11111_111110_11111;
    timing7[12][0] = 16'b11111_111110_11111;
    timing7[12][1] = 16'b00000_000000_00000;
    timing7[12][2] = 16'b00000_000000_00000;
    timing7[12][3] = 16'b11111_101110_00000;
    timing7[12][4] = 16'b11111_101110_00000;
    timing7[12][5] = 16'b11001_100100_00000;
    timing7[12][6] = 16'b11001_100100_00000;
    timing7[12][7] = 16'b11001_100100_00000;
    timing7[12][8] = 16'b11001_100100_00000;
    timing7[12][9] = 16'b11001_100100_00000;
    timing7[12][10] = 16'b11111_101110_00000;
    timing7[12][11] = 16'b11111_101110_00000;
    timing7[12][12] = 16'b00000_000000_00000;
    timing7[12][13] = 16'b00000_000000_00000;
    timing7[12][14] = 16'b11111_111110_11111;
    timing7[13][0] = 16'b11111_111110_11111;
    timing7[13][1] = 16'b00000_000000_00000;
    timing7[13][2] = 16'b00000_000000_00000;
    timing7[13][3] = 16'b00000_000000_00000;
    timing7[13][4] = 16'b00000_000000_00000;
    timing7[13][5] = 16'b11111_101110_00000;
    timing7[13][6] = 16'b11111_101110_00000;
    timing7[13][7] = 16'b11111_101110_00000;
    timing7[13][8] = 16'b11111_101110_00000;
    timing7[13][9] = 16'b11111_101110_00000;
    timing7[13][10] = 16'b00000_000000_00000;
    timing7[13][11] = 16'b00000_000000_00000;
    timing7[13][12] = 16'b00000_000000_00000;
    timing7[13][13] = 16'b00000_000000_00000;
    timing7[13][14] = 16'b11111_111110_11111;
    timing7[14][0] = 16'b11111_111110_11111;
    timing7[14][1] = 16'b11111_111110_11111;
    timing7[14][2] = 16'b11111_111110_11111;
    timing7[14][3] = 16'b11111_111110_11111;
    timing7[14][4] = 16'b11111_111110_11111;
    timing7[14][5] = 16'b11111_111110_11111;
    timing7[14][6] = 16'b11111_111110_11111;
    timing7[14][7] = 16'b11111_111110_11111;
    timing7[14][8] = 16'b11111_111110_11111;
    timing7[14][9] = 16'b11111_111110_11111;
    timing7[14][10] = 16'b11111_111110_11111;
    timing7[14][11] = 16'b11111_111110_11111;
    timing7[14][12] = 16'b11111_111110_11111;
    timing7[14][13] = 16'b11111_111110_11111;
    timing7[14][14] = 16'b11111_111110_11111;
    
    timing8[0][0] = 16'b11111_111110_11111;
    timing8[0][1] = 16'b11111_111110_11111;
    timing8[0][2] = 16'b11111_111110_11111;
    timing8[0][3] = 16'b11111_111110_11111;
    timing8[0][4] = 16'b11111_111110_11111;
    timing8[0][5] = 16'b11111_111110_11111;
    timing8[0][6] = 16'b11111_111110_11111;
    timing8[0][7] = 16'b11111_111110_11111;
    timing8[0][8] = 16'b11111_111110_11111;
    timing8[0][9] = 16'b11111_111110_11111;
    timing8[0][10] = 16'b11111_111110_11111;
    timing8[0][11] = 16'b11111_111110_11111;
    timing8[0][12] = 16'b11111_111110_11111;
    timing8[0][13] = 16'b11111_111110_11111;
    timing8[0][14] = 16'b11111_111110_11111;
    timing8[1][0] = 16'b11111_111110_11111;
    timing8[1][1] = 16'b00000_000000_00000;
    timing8[1][2] = 16'b00000_000000_00000;
    timing8[1][3] = 16'b00000_000000_00000;
    timing8[1][4] = 16'b00000_000000_00000;
    timing8[1][5] = 16'b11111_101110_00000;
    timing8[1][6] = 16'b11111_101110_00000;
    timing8[1][7] = 16'b11111_101110_00000;
    timing8[1][8] = 16'b11111_101110_00000;
    timing8[1][9] = 16'b11111_101110_00000;
    timing8[1][10] = 16'b00000_000000_00000;
    timing8[1][11] = 16'b00000_000000_00000;
    timing8[1][12] = 16'b00000_000000_00000;
    timing8[1][13] = 16'b00000_000000_00000;
    timing8[1][14] = 16'b11111_111110_11111;
    timing8[2][0] = 16'b11111_111110_11111;
    timing8[2][1] = 16'b00000_000000_00000;
    timing8[2][2] = 16'b00000_000000_00000;
    timing8[2][3] = 16'b11111_101110_00000;
    timing8[2][4] = 16'b11111_101110_00000;
    timing8[2][5] = 16'b11001_100100_00000;
    timing8[2][6] = 16'b11001_100100_00000;
    timing8[2][7] = 16'b11001_100100_00000;
    timing8[2][8] = 16'b11001_100100_00000;
    timing8[2][9] = 16'b11001_100100_00000;
    timing8[2][10] = 16'b11111_101110_00000;
    timing8[2][11] = 16'b11111_101110_00000;
    timing8[2][12] = 16'b00000_000000_00000;
    timing8[2][13] = 16'b00000_000000_00000;
    timing8[2][14] = 16'b11111_111110_11111;
    timing8[3][0] = 16'b11111_111110_11111;
    timing8[3][1] = 16'b00000_000000_00000;
    timing8[3][2] = 16'b11111_101110_00000;
    timing8[3][3] = 16'b11111_101110_00000;
    timing8[3][4] = 16'b11001_100100_00000;
    timing8[3][5] = 16'b11111_111110_11111;
    timing8[3][6] = 16'b11111_111110_11111;
    timing8[3][7] = 16'b11111_111110_11111;
    timing8[3][8] = 16'b11111_111110_11111;
    timing8[3][9] = 16'b11111_111110_11111;
    timing8[3][10] = 16'b11001_100100_00000;
    timing8[3][11] = 16'b11111_101110_00000;
    timing8[3][12] = 16'b11111_101110_00000;
    timing8[3][13] = 16'b00000_000000_00000;
    timing8[3][14] = 16'b11111_111110_11111;
    timing8[4][0] = 16'b11111_111110_11111;
    timing8[4][1] = 16'b00000_000000_00000;
    timing8[4][2] = 16'b11111_101110_00000;
    timing8[4][3] = 16'b11001_100100_00000;
    timing8[4][4] = 16'b11111_111110_11111;
    timing8[4][5] = 16'b00111_001111_00111;
    timing8[4][6] = 16'b11111_111110_11111;
    timing8[4][7] = 16'b11111_111110_11111;
    timing8[4][8] = 16'b11111_111110_11111;
    timing8[4][9] = 16'b11111_111110_11111;
    timing8[4][10] = 16'b11111_111110_11111;
    timing8[4][11] = 16'b11001_100100_00000;
    timing8[4][12] = 16'b11111_101110_00000;
    timing8[4][13] = 16'b00000_000000_00000;
    timing8[4][14] = 16'b11111_111110_11111;
    timing8[5][0] = 16'b11111_111110_11111;
    timing8[5][1] = 16'b11111_101110_00000;
    timing8[5][2] = 16'b11001_100100_00000;
    timing8[5][3] = 16'b11111_111110_11111;
    timing8[5][4] = 16'b11111_111110_11111;
    timing8[5][5] = 16'b00111_001111_00111;
    timing8[5][6] = 16'b11111_111110_11111;
    timing8[5][7] = 16'b11111_111110_11111;
    timing8[5][8] = 16'b11111_111110_11111;
    timing8[5][9] = 16'b11111_111110_11111;
    timing8[5][10] = 16'b11111_111110_11111;
    timing8[5][11] = 16'b11111_111110_11111;
    timing8[5][12] = 16'b11001_100100_00000;
    timing8[5][13] = 16'b11111_101110_00000;
    timing8[5][14] = 16'b11111_111110_11111;
    timing8[6][0] = 16'b11111_111110_11111;
    timing8[6][1] = 16'b11111_101110_00000;
    timing8[6][2] = 16'b11001_100100_00000;
    timing8[6][3] = 16'b11111_111110_11111;
    timing8[6][4] = 16'b11111_111110_11111;
    timing8[6][5] = 16'b11111_111110_11111;
    timing8[6][6] = 16'b00111_001111_00111;
    timing8[6][7] = 16'b11111_111110_11111;
    timing8[6][8] = 16'b11111_111110_11111;
    timing8[6][9] = 16'b11111_111110_11111;
    timing8[6][10] = 16'b11111_111110_11111;
    timing8[6][11] = 16'b11111_111110_11111;
    timing8[6][12] = 16'b11001_100100_00000;
    timing8[6][13] = 16'b11111_101110_00000;
    timing8[6][14] = 16'b11111_111110_11111;
    timing8[7][0] = 16'b11111_111110_11111;
    timing8[7][1] = 16'b11111_101110_00000;
    timing8[7][2] = 16'b11001_100100_00000;
    timing8[7][3] = 16'b11111_111110_11111;
    timing8[7][4] = 16'b11111_111110_11111;
    timing8[7][5] = 16'b11111_111110_11111;
    timing8[7][6] = 16'b11111_111110_11111;
    timing8[7][7] = 16'b00000_000000_00000;
    timing8[7][8] = 16'b00000_000000_00000;
    timing8[7][9] = 16'b00000_000000_00000;
    timing8[7][10] = 16'b00000_000000_00000;
    timing8[7][11] = 16'b11111_111110_11111;
    timing8[7][12] = 16'b11001_100100_00000;
    timing8[7][13] = 16'b11111_101110_00000;
    timing8[7][14] = 16'b11111_111110_11111;
    timing8[8][0] = 16'b11111_111110_11111;
    timing8[8][1] = 16'b11111_101110_00000;
    timing8[8][2] = 16'b11001_100100_00000;
    timing8[8][3] = 16'b11111_111110_11111;
    timing8[8][4] = 16'b11111_111110_11111;
    timing8[8][5] = 16'b11111_111110_11111;
    timing8[8][6] = 16'b11111_111110_11111;
    timing8[8][7] = 16'b11111_111110_11111;
    timing8[8][8] = 16'b11111_111110_11111;
    timing8[8][9] = 16'b11111_111110_11111;
    timing8[8][10] = 16'b11111_111110_11111;
    timing8[8][11] = 16'b11111_111110_11111;
    timing8[8][12] = 16'b11001_100100_00000;
    timing8[8][13] = 16'b11111_101110_00000;
    timing8[8][14] = 16'b11111_111110_11111;
    timing8[9][0] = 16'b11111_111110_11111;
    timing8[9][1] = 16'b11111_101110_00000;
    timing8[9][2] = 16'b11001_100100_00000;
    timing8[9][3] = 16'b11111_111110_11111;
    timing8[9][4] = 16'b11111_111110_11111;
    timing8[9][5] = 16'b11111_111110_11111;
    timing8[9][6] = 16'b11111_111110_11111;
    timing8[9][7] = 16'b11111_111110_11111;
    timing8[9][8] = 16'b11111_111110_11111;
    timing8[9][9] = 16'b11111_111110_11111;
    timing8[9][10] = 16'b11111_111110_11111;
    timing8[9][11] = 16'b11111_111110_11111;
    timing8[9][12] = 16'b11001_100100_00000;
    timing8[9][13] = 16'b11111_101110_00000;
    timing8[9][14] = 16'b11111_111110_11111;
    timing8[10][0] = 16'b11111_111110_11111;
    timing8[10][1] = 16'b00000_000000_00000;
    timing8[10][2] = 16'b11111_101110_00000;
    timing8[10][3] = 16'b11001_100100_00000;
    timing8[10][4] = 16'b11111_111110_11111;
    timing8[10][5] = 16'b11111_111110_11111;
    timing8[10][6] = 16'b11111_111110_11111;
    timing8[10][7] = 16'b11111_111110_11111;
    timing8[10][8] = 16'b11111_111110_11111;
    timing8[10][9] = 16'b11111_111110_11111;
    timing8[10][10] = 16'b11111_111110_11111;
    timing8[10][11] = 16'b11001_100100_00000;
    timing8[10][12] = 16'b11111_101110_00000;
    timing8[10][13] = 16'b00000_000000_00000;
    timing8[10][14] = 16'b11111_111110_11111;
    timing8[11][0] = 16'b11111_111110_11111;
    timing8[11][1] = 16'b00000_000000_00000;
    timing8[11][2] = 16'b11111_101110_00000;
    timing8[11][3] = 16'b11111_101110_00000;
    timing8[11][4] = 16'b11001_100100_00000;
    timing8[11][5] = 16'b11111_111110_11111;
    timing8[11][6] = 16'b11111_111110_11111;
    timing8[11][7] = 16'b11111_111110_11111;
    timing8[11][8] = 16'b11111_111110_11111;
    timing8[11][9] = 16'b11111_111110_11111;
    timing8[11][10] = 16'b11001_100100_00000;
    timing8[11][11] = 16'b11111_101110_00000;
    timing8[11][12] = 16'b11111_101110_00000;
    timing8[11][13] = 16'b00000_000000_00000;
    timing8[11][14] = 16'b11111_111110_11111;
    timing8[12][0] = 16'b11111_111110_11111;
    timing8[12][1] = 16'b00000_000000_00000;
    timing8[12][2] = 16'b00000_000000_00000;
    timing8[12][3] = 16'b11111_101110_00000;
    timing8[12][4] = 16'b11111_101110_00000;
    timing8[12][5] = 16'b11001_100100_00000;
    timing8[12][6] = 16'b11001_100100_00000;
    timing8[12][7] = 16'b11001_100100_00000;
    timing8[12][8] = 16'b11001_100100_00000;
    timing8[12][9] = 16'b11001_100100_00000;
    timing8[12][10] = 16'b11111_101110_00000;
    timing8[12][11] = 16'b11111_101110_00000;
    timing8[12][12] = 16'b00000_000000_00000;
    timing8[12][13] = 16'b00000_000000_00000;
    timing8[12][14] = 16'b11111_111110_11111;
    timing8[13][0] = 16'b11111_111110_11111;
    timing8[13][1] = 16'b00000_000000_00000;
    timing8[13][2] = 16'b00000_000000_00000;
    timing8[13][3] = 16'b00000_000000_00000;
    timing8[13][4] = 16'b00000_000000_00000;
    timing8[13][5] = 16'b11111_101110_00000;
    timing8[13][6] = 16'b11111_101110_00000;
    timing8[13][7] = 16'b11111_101110_00000;
    timing8[13][8] = 16'b11111_101110_00000;
    timing8[13][9] = 16'b11111_101110_00000;
    timing8[13][10] = 16'b00000_000000_00000;
    timing8[13][11] = 16'b00000_000000_00000;
    timing8[13][12] = 16'b00000_000000_00000;
    timing8[13][13] = 16'b00000_000000_00000;
    timing8[13][14] = 16'b11111_111110_11111;
    timing8[14][0] = 16'b11111_111110_11111;
    timing8[14][1] = 16'b11111_111110_11111;
    timing8[14][2] = 16'b11111_111110_11111;
    timing8[14][3] = 16'b11111_111110_11111;
    timing8[14][4] = 16'b11111_111110_11111;
    timing8[14][5] = 16'b11111_111110_11111;
    timing8[14][6] = 16'b11111_111110_11111;
    timing8[14][7] = 16'b11111_111110_11111;
    timing8[14][8] = 16'b11111_111110_11111;
    timing8[14][9] = 16'b11111_111110_11111;
    timing8[14][10] = 16'b11111_111110_11111;
    timing8[14][11] = 16'b11111_111110_11111;
    timing8[14][12] = 16'b11111_111110_11111;
    timing8[14][13] = 16'b11111_111110_11111;
    timing8[14][14] = 16'b11111_111110_11111;
    
    
    // FHKJSDFK
    timing9[0][0] = 16'b11111_111110_11111;
    timing9[0][1] = 16'b11111_111110_11111;
    timing9[0][2] = 16'b11111_111110_11111;
    timing9[0][3] = 16'b11111_111110_11111;
    timing9[0][4] = 16'b11111_111110_11111;
    timing9[0][5] = 16'b11111_111110_11111;
    timing9[0][6] = 16'b11111_111110_11111;
    timing9[0][7] = 16'b11111_111110_11111;
    timing9[0][8] = 16'b11111_111110_11111;
    timing9[0][9] = 16'b11111_111110_11111;
    timing9[0][10] = 16'b11111_111110_11111;
    timing9[0][11] = 16'b11111_111110_11111;
    timing9[0][12] = 16'b11111_111110_11111;
    timing9[0][13] = 16'b11111_111110_11111;
    timing9[0][14] = 16'b11111_111110_11111;
    timing9[1][0] = 16'b11111_111110_11111;
    timing9[1][1] = 16'b00000_000000_00000;
    timing9[1][2] = 16'b00000_000000_00000;
    timing9[1][3] = 16'b00000_000000_00000;
    timing9[1][4] = 16'b00000_000000_00000;
    timing9[1][5] = 16'b11111_101110_00000;
    timing9[1][6] = 16'b11111_101110_00000;
    timing9[1][7] = 16'b11111_101110_00000;
    timing9[1][8] = 16'b11111_101110_00000;
    timing9[1][9] = 16'b11111_101110_00000;
    timing9[1][10] = 16'b00000_000000_00000;
    timing9[1][11] = 16'b00000_000000_00000;
    timing9[1][12] = 16'b00000_000000_00000;
    timing9[1][13] = 16'b00000_000000_00000;
    timing9[1][14] = 16'b11111_111110_11111;
    timing9[2][0] = 16'b11111_111110_11111;
    timing9[2][1] = 16'b00000_000000_00000;
    timing9[2][2] = 16'b00000_000000_00000;
    timing9[2][3] = 16'b11111_101110_00000;
    timing9[2][4] = 16'b11111_101110_00000;
    timing9[2][5] = 16'b11001_100100_00000;
    timing9[2][6] = 16'b11001_100100_00000;
    timing9[2][7] = 16'b11001_100100_00000;
    timing9[2][8] = 16'b11001_100100_00000;
    timing9[2][9] = 16'b11001_100100_00000;
    timing9[2][10] = 16'b11111_101110_00000;
    timing9[2][11] = 16'b11111_101110_00000;
    timing9[2][12] = 16'b00000_000000_00000;
    timing9[2][13] = 16'b00000_000000_00000;
    timing9[2][14] = 16'b11111_111110_11111;
    timing9[3][0] = 16'b11111_111110_11111;
    timing9[3][1] = 16'b00000_000000_00000;
    timing9[3][2] = 16'b11111_101110_00000;
    timing9[3][3] = 16'b11111_101110_00000;
    timing9[3][4] = 16'b11001_100100_00000;
    timing9[3][5] = 16'b11111_111110_11111;
    timing9[3][6] = 16'b11111_111110_11111;
    timing9[3][7] = 16'b00111_001111_00111;
    timing9[3][8] = 16'b11111_111110_11111;
    timing9[3][9] = 16'b11111_111110_11111;
    timing9[3][10] = 16'b11001_100100_00000;
    timing9[3][11] = 16'b11111_101110_00000;
    timing9[3][12] = 16'b11111_101110_00000;
    timing9[3][13] = 16'b00000_000000_00000;
    timing9[3][14] = 16'b11111_111110_11111;
    timing9[4][0] = 16'b11111_111110_11111;
    timing9[4][1] = 16'b00000_000000_00000;
    timing9[4][2] = 16'b11111_101110_00000;
    timing9[4][3] = 16'b11001_100100_00000;
    timing9[4][4] = 16'b11111_111110_11111;
    timing9[4][5] = 16'b11111_111110_11111;
    timing9[4][6] = 16'b11111_111110_11111;
    timing9[4][7] = 16'b00111_001111_00111;
    timing9[4][8] = 16'b11111_111110_11111;
    timing9[4][9] = 16'b11111_111110_11111;
    timing9[4][10] = 16'b11111_111110_11111;
    timing9[4][11] = 16'b11001_100100_00000;
    timing9[4][12] = 16'b11111_101110_00000;
    timing9[4][13] = 16'b00000_000000_00000;
    timing9[4][14] = 16'b11111_111110_11111;
    timing9[5][0] = 16'b11111_111110_11111;
    timing9[5][1] = 16'b11111_101110_00000;
    timing9[5][2] = 16'b11001_100100_00000;
    timing9[5][3] = 16'b11111_111110_11111;
    timing9[5][4] = 16'b11111_111110_11111;
    timing9[5][5] = 16'b11111_111110_11111;
    timing9[5][6] = 16'b11111_111110_11111;
    timing9[5][7] = 16'b00111_001111_00111;
    timing9[5][8] = 16'b11111_111110_11111;
    timing9[5][9] = 16'b11111_111110_11111;
    timing9[5][10] = 16'b11111_111110_11111;
    timing9[5][11] = 16'b11111_111110_11111;
    timing9[5][12] = 16'b11001_100100_00000;
    timing9[5][13] = 16'b11111_101110_00000;
    timing9[5][14] = 16'b11111_111110_11111;
    timing9[6][0] = 16'b11111_111110_11111;
    timing9[6][1] = 16'b11111_101110_00000;
    timing9[6][2] = 16'b11001_100100_00000;
    timing9[6][3] = 16'b11111_111110_11111;
    timing9[6][4] = 16'b11111_111110_11111;
    timing9[6][5] = 16'b11111_111110_11111;
    timing9[6][6] = 16'b11111_111110_11111;
    timing9[6][7] = 16'b00111_001111_00111;
    timing9[6][8] = 16'b11111_111110_11111;
    timing9[6][9] = 16'b11111_111110_11111;
    timing9[6][10] = 16'b11111_111110_11111;
    timing9[6][11] = 16'b11111_111110_11111;
    timing9[6][12] = 16'b11001_100100_00000;
    timing9[6][13] = 16'b11111_101110_00000;
    timing9[6][14] = 16'b11111_111110_11111;
    timing9[7][0] = 16'b11111_111110_11111;
    timing9[7][1] = 16'b11111_101110_00000;
    timing9[7][2] = 16'b11001_100100_00000;
    timing9[7][3] = 16'b11111_111110_11111;
    timing9[7][4] = 16'b11111_111110_11111;
    timing9[7][5] = 16'b11111_111110_11111;
    timing9[7][6] = 16'b11111_111110_11111;
    timing9[7][7] = 16'b00000_000000_00000;
    timing9[7][8] = 16'b00000_000000_00000;
    timing9[7][9] = 16'b00000_000000_00000;
    timing9[7][10] = 16'b00000_000000_00000;
    timing9[7][11] = 16'b11111_111110_11111;
    timing9[7][12] = 16'b11001_100100_00000;
    timing9[7][13] = 16'b11111_101110_00000;
    timing9[7][14] = 16'b11111_111110_11111;
    timing9[8][0] = 16'b11111_111110_11111;
    timing9[8][1] = 16'b11111_101110_00000;
    timing9[8][2] = 16'b11001_100100_00000;
    timing9[8][3] = 16'b11111_111110_11111;
    timing9[8][4] = 16'b11111_111110_11111;
    timing9[8][5] = 16'b11111_111110_11111;
    timing9[8][6] = 16'b11111_111110_11111;
    timing9[8][7] = 16'b11111_111110_11111;
    timing9[8][8] = 16'b11111_111110_11111;
    timing9[8][9] = 16'b11111_111110_11111;
    timing9[8][10] = 16'b11111_111110_11111;
    timing9[8][11] = 16'b11111_111110_11111;
    timing9[8][12] = 16'b11001_100100_00000;
    timing9[8][13] = 16'b11111_101110_00000;
    timing9[8][14] = 16'b11111_111110_11111;
    timing9[9][0] = 16'b11111_111110_11111;
    timing9[9][1] = 16'b11111_101110_00000;
    timing9[9][2] = 16'b11001_100100_00000;
    timing9[9][3] = 16'b11111_111110_11111;
    timing9[9][4] = 16'b11111_111110_11111;
    timing9[9][5] = 16'b11111_111110_11111;
    timing9[9][6] = 16'b11111_111110_11111;
    timing9[9][7] = 16'b11111_111110_11111;
    timing9[9][8] = 16'b11111_111110_11111;
    timing9[9][9] = 16'b11111_111110_11111;
    timing9[9][10] = 16'b11111_111110_11111;
    timing9[9][11] = 16'b11111_111110_11111;
    timing9[9][12] = 16'b11001_100100_00000;
    timing9[9][13] = 16'b11111_101110_00000;
    timing9[9][14] = 16'b11111_111110_11111;
    timing9[10][0] = 16'b11111_111110_11111;
    timing9[10][1] = 16'b00000_000000_00000;
    timing9[10][2] = 16'b11111_101110_00000;
    timing9[10][3] = 16'b11001_100100_00000;
    timing9[10][4] = 16'b11111_111110_11111;
    timing9[10][5] = 16'b11111_111110_11111;
    timing9[10][6] = 16'b11111_111110_11111;
    timing9[10][7] = 16'b11111_111110_11111;
    timing9[10][8] = 16'b11111_111110_11111;
    timing9[10][9] = 16'b11111_111110_11111;
    timing9[10][10] = 16'b11111_111110_11111;
    timing9[10][11] = 16'b11001_100100_00000;
    timing9[10][12] = 16'b11111_101110_00000;
    timing9[10][13] = 16'b00000_000000_00000;
    timing9[10][14] = 16'b11111_111110_11111;
    timing9[11][0] = 16'b11111_111110_11111;
    timing9[11][1] = 16'b00000_000000_00000;
    timing9[11][2] = 16'b11111_101110_00000;
    timing9[11][3] = 16'b11111_101110_00000;
    timing9[11][4] = 16'b11001_100100_00000;
    timing9[11][5] = 16'b11111_111110_11111;
    timing9[11][6] = 16'b11111_111110_11111;
    timing9[11][7] = 16'b11111_111110_11111;
    timing9[11][8] = 16'b11111_111110_11111;
    timing9[11][9] = 16'b11111_111110_11111;
    timing9[11][10] = 16'b11001_100100_00000;
    timing9[11][11] = 16'b11111_101110_00000;
    timing9[11][12] = 16'b11111_101110_00000;
    timing9[11][13] = 16'b00000_000000_00000;
    timing9[11][14] = 16'b11111_111110_11111;
    timing9[12][0] = 16'b11111_111110_11111;
    timing9[12][1] = 16'b00000_000000_00000;
    timing9[12][2] = 16'b00000_000000_00000;
    timing9[12][3] = 16'b11111_101110_00000;
    timing9[12][4] = 16'b11111_101110_00000;
    timing9[12][5] = 16'b11001_100100_00000;
    timing9[12][6] = 16'b11001_100100_00000;
    timing9[12][7] = 16'b11001_100100_00000;
    timing9[12][8] = 16'b11001_100100_00000;
    timing9[12][9] = 16'b11001_100100_00000;
    timing9[12][10] = 16'b11111_101110_00000;
    timing9[12][11] = 16'b11111_101110_00000;
    timing9[12][12] = 16'b00000_000000_00000;
    timing9[12][13] = 16'b00000_000000_00000;
    timing9[12][14] = 16'b11111_111110_11111;
    timing9[13][0] = 16'b11111_111110_11111;
    timing9[13][1] = 16'b00000_000000_00000;
    timing9[13][2] = 16'b00000_000000_00000;
    timing9[13][3] = 16'b00000_000000_00000;
    timing9[13][4] = 16'b00000_000000_00000;
    timing9[13][5] = 16'b11111_101110_00000;
    timing9[13][6] = 16'b11111_101110_00000;
    timing9[13][7] = 16'b11111_101110_00000;
    timing9[13][8] = 16'b11111_101110_00000;
    timing9[13][9] = 16'b11111_101110_00000;
    timing9[13][10] = 16'b00000_000000_00000;
    timing9[13][11] = 16'b00000_000000_00000;
    timing9[13][12] = 16'b00000_000000_00000;
    timing9[13][13] = 16'b00000_000000_00000;
    timing9[13][14] = 16'b11111_111110_11111;
    timing9[14][0] = 16'b11111_111110_11111;
    timing9[14][1] = 16'b11111_111110_11111;
    timing9[14][2] = 16'b11111_111110_11111;
    timing9[14][3] = 16'b11111_111110_11111;
    timing9[14][4] = 16'b11111_111110_11111;
    timing9[14][5] = 16'b11111_111110_11111;
    timing9[14][6] = 16'b11111_111110_11111;
    timing9[14][7] = 16'b11111_111110_11111;
    timing9[14][8] = 16'b11111_111110_11111;
    timing9[14][9] = 16'b11111_111110_11111;
    timing9[14][10] = 16'b11111_111110_11111;
    timing9[14][11] = 16'b11111_111110_11111;
    timing9[14][12] = 16'b11111_111110_11111;
    timing9[14][13] = 16'b11111_111110_11111;
    timing9[14][14] = 16'b11111_111110_11111;
    
    chop_empty[0][0] = 16'b11111_111110_11111;
    chop_empty[0][1] = 16'b11111_111110_11111;
    chop_empty[0][2] = 16'b11111_111110_11111;
    chop_empty[0][3] = 16'b11111_111110_11111;
    chop_empty[0][4] = 16'b11111_111110_11111;
    chop_empty[0][5] = 16'b11111_111110_11111;
    chop_empty[0][6] = 16'b11111_111110_11111;
    chop_empty[0][7] = 16'b11111_111110_11111;
    chop_empty[0][8] = 16'b11111_111110_11111;
    chop_empty[0][9] = 16'b11111_111110_11111;
    chop_empty[0][10] = 16'b11111_111110_11111;
    chop_empty[0][11] = 16'b11111_111110_11111;
    chop_empty[0][12] = 16'b11111_111110_11111;
    chop_empty[0][13] = 16'b11111_111110_11111;
    chop_empty[0][14] = 16'b11111_111110_11111;
    chop_empty[1][0] = 16'b11111_111110_11111;
    chop_empty[1][1] = 16'b00000_000000_00000;
    chop_empty[1][2] = 16'b00000_000000_00000;
    chop_empty[1][3] = 16'b00000_000000_00000;
    chop_empty[1][4] = 16'b00000_000000_00000;
    chop_empty[1][5] = 16'b00000_000000_00000;
    chop_empty[1][6] = 16'b00000_000000_00000;
    chop_empty[1][7] = 16'b00000_000000_00000;
    chop_empty[1][8] = 16'b00000_000000_00000;
    chop_empty[1][9] = 16'b00000_000000_00000;
    chop_empty[1][10] = 16'b00000_000000_00000;
    chop_empty[1][11] = 16'b00000_000000_00000;
    chop_empty[1][12] = 16'b00000_000000_00000;
    chop_empty[1][13] = 16'b00000_000000_00000;
    chop_empty[1][14] = 16'b11111_111110_11111;
    chop_empty[2][0] = 16'b11111_111110_11111;
    chop_empty[2][1] = 16'b00000_000000_00000;
    chop_empty[2][2] = 16'b00000_000000_00000;
    chop_empty[2][3] = 16'b00000_000000_00000;
    chop_empty[2][4] = 16'b00000_000000_00000;
    chop_empty[2][5] = 16'b00000_000000_00000;
    chop_empty[2][6] = 16'b00000_000000_00000;
    chop_empty[2][7] = 16'b00000_000000_00000;
    chop_empty[2][8] = 16'b00000_000000_00000;
    chop_empty[2][9] = 16'b00000_000000_00000;
    chop_empty[2][10] = 16'b00000_000000_00000;
    chop_empty[2][11] = 16'b00000_000000_00000;
    chop_empty[2][12] = 16'b00000_000000_00000;
    chop_empty[2][13] = 16'b00000_000000_00000;
    chop_empty[2][14] = 16'b11111_111110_11111;
    chop_empty[3][0] = 16'b11111_111110_11111;
    chop_empty[3][1] = 16'b00000_000000_00000;
    chop_empty[3][2] = 16'b11111_110011_01110;
    chop_empty[3][3] = 16'b11111_110011_01110;
    chop_empty[3][4] = 16'b11111_110011_01110;
    chop_empty[3][5] = 16'b11111_110011_01110;
    chop_empty[3][6] = 16'b11111_110011_01110;
    chop_empty[3][7] = 16'b11111_110011_01110;
    chop_empty[3][8] = 16'b11111_110011_01110;
    chop_empty[3][9] = 16'b11111_110011_01110;
    chop_empty[3][10] = 16'b11111_110011_01110;
    chop_empty[3][11] = 16'b11111_110011_01110;
    chop_empty[3][12] = 16'b11111_110011_01110;
    chop_empty[3][13] = 16'b00000_000000_00000;
    chop_empty[3][14] = 16'b11111_111110_11111;
    chop_empty[4][0] = 16'b11111_111110_11111;
    chop_empty[4][1] = 16'b00000_000000_00000;
    chop_empty[4][2] = 16'b11111_110011_01110;
    chop_empty[4][3] = 16'b11111_110011_01110;
    chop_empty[4][4] = 16'b11111_110011_01110;
    chop_empty[4][5] = 16'b11111_110011_01110;
    chop_empty[4][6] = 16'b11111_110011_01110;
    chop_empty[4][7] = 16'b11111_110011_01110;
    chop_empty[4][8] = 16'b11111_110011_01110;
    chop_empty[4][9] = 16'b11111_110011_01110;
    chop_empty[4][10] = 16'b11111_110011_01110;
    chop_empty[4][11] = 16'b11111_110011_01110;
    chop_empty[4][12] = 16'b11111_110011_01110;
    chop_empty[4][13] = 16'b00000_000000_00000;
    chop_empty[4][14] = 16'b11111_111110_11111;
    chop_empty[5][0] = 16'b11111_111110_11111;
    chop_empty[5][1] = 16'b00000_000000_00000;
    chop_empty[5][2] = 16'b11111_110011_01110;
    chop_empty[5][3] = 16'b11111_110011_01110;
    chop_empty[5][4] = 16'b11111_110011_01110;
    chop_empty[5][5] = 16'b11111_110011_01110;
    chop_empty[5][6] = 16'b11111_110011_01110;
    chop_empty[5][7] = 16'b11111_110011_01110;
    chop_empty[5][8] = 16'b11111_110011_01110;
    chop_empty[5][9] = 16'b11111_110011_01110;
    chop_empty[5][10] = 16'b11111_110011_01110;
    chop_empty[5][11] = 16'b11111_110011_01110;
    chop_empty[5][12] = 16'b11111_110011_01110;
    chop_empty[5][13] = 16'b00000_000000_00000;
    chop_empty[5][14] = 16'b11111_111110_11111;
    chop_empty[6][0] = 16'b11111_111110_11111;
    chop_empty[6][1] = 16'b00000_000000_00000;
    chop_empty[6][2] = 16'b11111_110011_01110;
    chop_empty[6][3] = 16'b11111_110011_01110;
    chop_empty[6][4] = 16'b11111_110011_01110;
    chop_empty[6][5] = 16'b11111_110011_01110;
    chop_empty[6][6] = 16'b11111_110011_01110;
    chop_empty[6][7] = 16'b11111_110011_01110;
    chop_empty[6][8] = 16'b11111_110011_01110;
    chop_empty[6][9] = 16'b11111_110011_01110;
    chop_empty[6][10] = 16'b11111_110011_01110;
    chop_empty[6][11] = 16'b11111_110011_01110;
    chop_empty[6][12] = 16'b11111_110011_01110;
    chop_empty[6][13] = 16'b00000_000000_00000;
    chop_empty[6][14] = 16'b11111_111110_11111;
    chop_empty[7][0] = 16'b11111_111110_11111;
    chop_empty[7][1] = 16'b00000_000000_00000;
    chop_empty[7][2] = 16'b11111_110011_01110;
    chop_empty[7][3] = 16'b11111_110011_01110;
    chop_empty[7][4] = 16'b11111_110011_01110;
    chop_empty[7][5] = 16'b11111_110011_01110;
    chop_empty[7][6] = 16'b11111_110011_01110;
    chop_empty[7][7] = 16'b11111_110011_01110;
    chop_empty[7][8] = 16'b11111_110011_01110;
    chop_empty[7][9] = 16'b11111_110011_01110;
    chop_empty[7][10] = 16'b11111_110011_01110;
    chop_empty[7][11] = 16'b11111_110011_01110;
    chop_empty[7][12] = 16'b11111_110011_01110;
    chop_empty[7][13] = 16'b00000_000000_00000;
    chop_empty[7][14] = 16'b11111_111110_11111;
    chop_empty[8][0] = 16'b11111_111110_11111;
    chop_empty[8][1] = 16'b00000_000000_00000;
    chop_empty[8][2] = 16'b11111_110011_01110;
    chop_empty[8][3] = 16'b11111_110011_01110;
    chop_empty[8][4] = 16'b11111_110011_01110;
    chop_empty[8][5] = 16'b11111_110011_01110;
    chop_empty[8][6] = 16'b11111_110011_01110;
    chop_empty[8][7] = 16'b11111_110011_01110;
    chop_empty[8][8] = 16'b11111_110011_01110;
    chop_empty[8][9] = 16'b11111_110011_01110;
    chop_empty[8][10] = 16'b11111_110011_01110;
    chop_empty[8][11] = 16'b11111_110011_01110;
    chop_empty[8][12] = 16'b11111_110011_01110;
    chop_empty[8][13] = 16'b00000_000000_00000;
    chop_empty[8][14] = 16'b11111_111110_11111;
    chop_empty[9][0] = 16'b11111_111110_11111;
    chop_empty[9][1] = 16'b00000_000000_00000;
    chop_empty[9][2] = 16'b11111_110011_01110;
    chop_empty[9][3] = 16'b11111_110011_01110;
    chop_empty[9][4] = 16'b11111_110011_01110;
    chop_empty[9][5] = 16'b11111_110011_01110;
    chop_empty[9][6] = 16'b11111_110011_01110;
    chop_empty[9][7] = 16'b11111_110011_01110;
    chop_empty[9][8] = 16'b11111_110011_01110;
    chop_empty[9][9] = 16'b11111_110011_01110;
    chop_empty[9][10] = 16'b11111_110011_01110;
    chop_empty[9][11] = 16'b11111_110011_01110;
    chop_empty[9][12] = 16'b11111_110011_01110;
    chop_empty[9][13] = 16'b00000_000000_00000;
    chop_empty[9][14] = 16'b11111_111110_11111;
    chop_empty[10][0] = 16'b11111_111110_11111;
    chop_empty[10][1] = 16'b00000_000000_00000;
    chop_empty[10][2] = 16'b11111_110011_01110;
    chop_empty[10][3] = 16'b11111_110011_01110;
    chop_empty[10][4] = 16'b11111_110011_01110;
    chop_empty[10][5] = 16'b11111_110011_01110;
    chop_empty[10][6] = 16'b11111_110011_01110;
    chop_empty[10][7] = 16'b11111_110011_01110;
    chop_empty[10][8] = 16'b11111_110011_01110;
    chop_empty[10][9] = 16'b11111_110011_01110;
    chop_empty[10][10] = 16'b11111_110011_01110;
    chop_empty[10][11] = 16'b11111_110011_01110;
    chop_empty[10][12] = 16'b11111_110011_01110;
    chop_empty[10][13] = 16'b00000_000000_00000;
    chop_empty[10][14] = 16'b11111_111110_11111;
    chop_empty[11][0] = 16'b11111_111110_11111;
    chop_empty[11][1] = 16'b00000_000000_00000;
    chop_empty[11][2] = 16'b00000_000000_00000;
    chop_empty[11][3] = 16'b00000_000000_00000;
    chop_empty[11][4] = 16'b00000_000000_00000;
    chop_empty[11][5] = 16'b00000_000000_00000;
    chop_empty[11][6] = 16'b00000_000000_00000;
    chop_empty[11][7] = 16'b00000_000000_00000;
    chop_empty[11][8] = 16'b00000_000000_00000;
    chop_empty[11][9] = 16'b00000_000000_00000;
    chop_empty[11][10] = 16'b00000_000000_00000;
    chop_empty[11][11] = 16'b00000_000000_00000;
    chop_empty[11][12] = 16'b00000_000000_00000;
    chop_empty[11][13] = 16'b00000_000000_00000;
    chop_empty[11][14] = 16'b11111_111110_11111;
    chop_empty[12][0] = 16'b11111_111110_11111;
    chop_empty[12][1] = 16'b00000_000000_00000;
    chop_empty[12][2] = 16'b00000_000000_00000;
    chop_empty[12][3] = 16'b00000_000000_00000;
    chop_empty[12][4] = 16'b00000_000000_00000;
    chop_empty[12][5] = 16'b00000_000000_00000;
    chop_empty[12][6] = 16'b00000_000000_00000;
    chop_empty[12][7] = 16'b00000_000000_00000;
    chop_empty[12][8] = 16'b00000_000000_00000;
    chop_empty[12][9] = 16'b00000_000000_00000;
    chop_empty[12][10] = 16'b00000_000000_00000;
    chop_empty[12][11] = 16'b00000_000000_00000;
    chop_empty[12][12] = 16'b00000_000000_00000;
    chop_empty[12][13] = 16'b00000_000000_00000;
    chop_empty[12][14] = 16'b11111_111110_11111;
    chop_empty[13][0] = 16'b11111_111110_11111;
    chop_empty[13][1] = 16'b00000_000000_00000;
    chop_empty[13][2] = 16'b00000_000000_00000;
    chop_empty[13][3] = 16'b00000_000000_00000;
    chop_empty[13][4] = 16'b00000_000000_00000;
    chop_empty[13][5] = 16'b00000_000000_00000;
    chop_empty[13][6] = 16'b00000_000000_00000;
    chop_empty[13][7] = 16'b00000_000000_00000;
    chop_empty[13][8] = 16'b00000_000000_00000;
    chop_empty[13][9] = 16'b00000_000000_00000;
    chop_empty[13][10] = 16'b00000_000000_00000;
    chop_empty[13][11] = 16'b00000_000000_00000;
    chop_empty[13][12] = 16'b00000_000000_00000;
    chop_empty[13][13] = 16'b00000_000000_00000;
    chop_empty[13][14] = 16'b11111_111110_11111;
    chop_empty[14][0] = 16'b11111_111110_11111;
    chop_empty[14][1] = 16'b11111_111110_11111;
    chop_empty[14][2] = 16'b11111_111110_11111;
    chop_empty[14][3] = 16'b11111_111110_11111;
    chop_empty[14][4] = 16'b11111_111110_11111;
    chop_empty[14][5] = 16'b11111_111110_11111;
    chop_empty[14][6] = 16'b11111_111110_11111;
    chop_empty[14][7] = 16'b11111_111110_11111;
    chop_empty[14][8] = 16'b11111_111110_11111;
    chop_empty[14][9] = 16'b11111_111110_11111;
    chop_empty[14][10] = 16'b11111_111110_11111;
    chop_empty[14][11] = 16'b11111_111110_11111;
    chop_empty[14][12] = 16'b11111_111110_11111;
    chop_empty[14][13] = 16'b11111_111110_11111;
    chop_empty[14][14] = 16'b11111_111110_11111;
    
    chop_full[0][0] = 16'b11111_111110_11111;
    chop_full[0][1] = 16'b11111_111110_11111;
    chop_full[0][2] = 16'b11111_111110_11111;
    chop_full[0][3] = 16'b11111_111110_11111;
    chop_full[0][4] = 16'b11111_111110_11111;
    chop_full[0][5] = 16'b11111_111110_11111;
    chop_full[0][6] = 16'b11111_111110_11111;
    chop_full[0][7] = 16'b11111_111110_11111;
    chop_full[0][8] = 16'b11111_111110_11111;
    chop_full[0][9] = 16'b11111_111110_11111;
    chop_full[0][10] = 16'b11111_111110_11111;
    chop_full[0][11] = 16'b11111_111110_11111;
    chop_full[0][12] = 16'b11111_111110_11111;
    chop_full[0][13] = 16'b11111_111110_11111;
    chop_full[0][14] = 16'b11111_111110_11111;
    chop_full[1][0] = 16'b11111_111110_11111;
    chop_full[1][1] = 16'b00000_000000_00000;
    chop_full[1][2] = 16'b00000_000000_00000;
    chop_full[1][3] = 16'b00000_000000_00000;
    chop_full[1][4] = 16'b00000_000000_00000;
    chop_full[1][5] = 16'b00000_000000_00000;
    chop_full[1][6] = 16'b00000_000000_00000;
    chop_full[1][7] = 16'b00000_000000_00000;
    chop_full[1][8] = 16'b00000_000000_00000;
    chop_full[1][9] = 16'b00000_000000_00000;
    chop_full[1][10] = 16'b00000_000000_00000;
    chop_full[1][11] = 16'b00000_000000_00000;
    chop_full[1][12] = 16'b00000_000000_00000;
    chop_full[1][13] = 16'b00000_000000_00000;
    chop_full[1][14] = 16'b11111_111110_11111;
    chop_full[2][0] = 16'b11111_111110_11111;
    chop_full[2][1] = 16'b00000_000000_00000;
    chop_full[2][2] = 16'b00000_000000_00000;
    chop_full[2][3] = 16'b00000_000000_00000;
    chop_full[2][4] = 16'b00000_000000_00000;
    chop_full[2][5] = 16'b00000_000000_00000;
    chop_full[2][6] = 16'b00000_000000_00000;
    chop_full[2][7] = 16'b00000_000000_00000;
    chop_full[2][8] = 16'b00000_000000_00000;
    chop_full[2][9] = 16'b00000_000000_00000;
    chop_full[2][10] = 16'b00000_000000_00000;
    chop_full[2][11] = 16'b00000_000000_00000;
    chop_full[2][12] = 16'b00000_000000_00000;
    chop_full[2][13] = 16'b00000_000000_00000;
    chop_full[2][14] = 16'b11111_111110_11111;
    chop_full[3][0] = 16'b11111_111110_11111;
    chop_full[3][1] = 16'b00000_000000_00000;
    chop_full[3][2] = 16'b11111_110011_01110;
    chop_full[3][3] = 16'b11111_110011_01110;
    chop_full[3][4] = 16'b11111_110011_01110;
    chop_full[3][5] = 16'b11111_110011_01110;
    chop_full[3][6] = 16'b11111_110011_01110;
    chop_full[3][7] = 16'b11111_110011_01110;
    chop_full[3][8] = 16'b11111_110011_01110;
    chop_full[3][9] = 16'b11111_110011_01110;
    chop_full[3][10] = 16'b11111_110011_01110;
    chop_full[3][11] = 16'b11111_110011_01110;
    chop_full[3][12] = 16'b11111_110011_01110;
    chop_full[3][13] = 16'b00000_000000_00000;
    chop_full[3][14] = 16'b11111_111110_11111;
    chop_full[4][0] = 16'b11111_111110_11111;
    chop_full[4][1] = 16'b00000_000000_00000;
    chop_full[4][2] = 16'b11111_110011_01110;
    chop_full[4][3] = 16'b11111_110011_01110;
    chop_full[4][4] = 16'b11111_110011_01110;
    chop_full[4][5] = 16'b10111_011111_00000;
    chop_full[4][6] = 16'b10111_011111_00000;
    chop_full[4][7] = 16'b10111_011111_00000;
    chop_full[4][8] = 16'b10111_011111_00000;
    chop_full[4][9] = 16'b10111_011111_00000;
    chop_full[4][10] = 16'b11111_110011_01110;
    chop_full[4][11] = 16'b11111_110011_01110;
    chop_full[4][12] = 16'b11111_110011_01110;
    chop_full[4][13] = 16'b00000_000000_00000;
    chop_full[4][14] = 16'b11111_111110_11111;
    chop_full[5][0] = 16'b11111_111110_11111;
    chop_full[5][1] = 16'b00000_000000_00000;
    chop_full[5][2] = 16'b11111_110011_01110;
    chop_full[5][3] = 16'b11111_110011_01110;
    chop_full[5][4] = 16'b10111_011111_00000;
    chop_full[5][5] = 16'b10111_011111_00000;
    chop_full[5][6] = 16'b10111_011111_00000;
    chop_full[5][7] = 16'b10111_011111_00000;
    chop_full[5][8] = 16'b10111_011111_00000;
    chop_full[5][9] = 16'b10111_011111_00000;
    chop_full[5][10] = 16'b10111_011111_00000;
    chop_full[5][11] = 16'b11111_110011_01110;
    chop_full[5][12] = 16'b11111_110011_01110;
    chop_full[5][13] = 16'b00000_000000_00000;
    chop_full[5][14] = 16'b11111_111110_11111;
    chop_full[6][0] = 16'b11111_111110_11111;
    chop_full[6][1] = 16'b00000_000000_00000;
    chop_full[6][2] = 16'b11111_110011_01110;
    chop_full[6][3] = 16'b10111_011111_00000;
    chop_full[6][4] = 16'b10111_011111_00000;
    chop_full[6][5] = 16'b10111_011111_00000;
    chop_full[6][6] = 16'b10111_011111_00000;
    chop_full[6][7] = 16'b10111_011111_00000;
    chop_full[6][8] = 16'b10111_011111_00000;
    chop_full[6][9] = 16'b10111_011111_00000;
    chop_full[6][10] = 16'b10111_011111_00000;
    chop_full[6][11] = 16'b10111_011111_00000;
    chop_full[6][12] = 16'b11111_110011_01110;
    chop_full[6][13] = 16'b00000_000000_00000;
    chop_full[6][14] = 16'b11111_111110_11111;
    chop_full[7][0] = 16'b11111_111110_11111;
    chop_full[7][1] = 16'b00000_000000_00000;
    chop_full[7][2] = 16'b11111_110011_01110;
    chop_full[7][3] = 16'b10111_011111_00000;
    chop_full[7][4] = 16'b10111_011111_00000;
    chop_full[7][5] = 16'b10111_011111_00000;
    chop_full[7][6] = 16'b10111_011111_00000;
    chop_full[7][7] = 16'b10111_011111_00000;
    chop_full[7][8] = 16'b10111_011111_00000;
    chop_full[7][9] = 16'b10111_011111_00000;
    chop_full[7][10] = 16'b10111_011111_00000;
    chop_full[7][11] = 16'b10111_011111_00000;
    chop_full[7][12] = 16'b11111_110011_01110;
    chop_full[7][13] = 16'b00000_000000_00000;
    chop_full[7][14] = 16'b11111_111110_11111;
    chop_full[8][0] = 16'b11111_111110_11111;
    chop_full[8][1] = 16'b00000_000000_00000;
    chop_full[8][2] = 16'b11111_110011_01110;
    chop_full[8][3] = 16'b10111_011111_00000;
    chop_full[8][4] = 16'b10111_011111_00000;
    chop_full[8][5] = 16'b10111_011111_00000;
    chop_full[8][6] = 16'b10111_011111_00000;
    chop_full[8][7] = 16'b10111_011111_00000;
    chop_full[8][8] = 16'b10111_011111_00000;
    chop_full[8][9] = 16'b10111_011111_00000;
    chop_full[8][10] = 16'b10111_011111_00000;
    chop_full[8][11] = 16'b10111_011111_00000;
    chop_full[8][12] = 16'b11111_110011_01110;
    chop_full[8][13] = 16'b00000_000000_00000;
    chop_full[8][14] = 16'b11111_111110_11111;
    chop_full[9][0] = 16'b11111_111110_11111;
    chop_full[9][1] = 16'b00000_000000_00000;
    chop_full[9][2] = 16'b11111_110011_01110;
    chop_full[9][3] = 16'b11111_110011_01110;
    chop_full[9][4] = 16'b10111_011111_00000;
    chop_full[9][5] = 16'b10111_011111_00000;
    chop_full[9][6] = 16'b10111_011111_00000;
    chop_full[9][7] = 16'b10111_011111_00000;
    chop_full[9][8] = 16'b10111_011111_00000;
    chop_full[9][9] = 16'b10111_011111_00000;
    chop_full[9][10] = 16'b10111_011111_00000;
    chop_full[9][11] = 16'b11111_110011_01110;
    chop_full[9][12] = 16'b11111_110011_01110;
    chop_full[9][13] = 16'b00000_000000_00000;
    chop_full[9][14] = 16'b11111_111110_11111;
    chop_full[10][0] = 16'b11111_111110_11111;
    chop_full[10][1] = 16'b00000_000000_00000;
    chop_full[10][2] = 16'b11111_110011_01110;
    chop_full[10][3] = 16'b11111_110011_01110;
    chop_full[10][4] = 16'b11111_110011_01110;
    chop_full[10][5] = 16'b10111_011111_00000;
    chop_full[10][6] = 16'b10111_011111_00000;
    chop_full[10][7] = 16'b10111_011111_00000;
    chop_full[10][8] = 16'b10111_011111_00000;
    chop_full[10][9] = 16'b10111_011111_00000;
    chop_full[10][10] = 16'b11111_110011_01110;
    chop_full[10][11] = 16'b11111_110011_01110;
    chop_full[10][12] = 16'b11111_110011_01110;
    chop_full[10][13] = 16'b00000_000000_00000;
    chop_full[10][14] = 16'b11111_111110_11111;
    chop_full[11][0] = 16'b11111_111110_11111;
    chop_full[11][1] = 16'b00000_000000_00000;
    chop_full[11][2] = 16'b11111_110011_01110;
    chop_full[11][3] = 16'b11111_110011_01110;
    chop_full[11][4] = 16'b11111_110011_01110;
    chop_full[11][5] = 16'b11111_110011_01110;
    chop_full[11][6] = 16'b11111_110011_01110;
    chop_full[11][7] = 16'b11111_110011_01110;
    chop_full[11][8] = 16'b11111_110011_01110;
    chop_full[11][9] = 16'b11111_110011_01110;
    chop_full[11][10] = 16'b11111_110011_01110;
    chop_full[11][11] = 16'b11111_110011_01110;
    chop_full[11][12] = 16'b11111_110011_01110;
    chop_full[11][13] = 16'b00000_000000_00000;
    chop_full[11][14] = 16'b11111_111110_11111;
    chop_full[12][0] = 16'b11111_111110_11111;
    chop_full[12][1] = 16'b00000_000000_00000;
    chop_full[12][2] = 16'b00000_000000_00000;
    chop_full[12][3] = 16'b00000_000000_00000;
    chop_full[12][4] = 16'b00000_000000_00000;
    chop_full[12][5] = 16'b00000_000000_00000;
    chop_full[12][6] = 16'b00000_000000_00000;
    chop_full[12][7] = 16'b00000_000000_00000;
    chop_full[12][8] = 16'b00000_000000_00000;
    chop_full[12][9] = 16'b00000_000000_00000;
    chop_full[12][10] = 16'b00000_000000_00000;
    chop_full[12][11] = 16'b00000_000000_00000;
    chop_full[12][12] = 16'b00000_000000_00000;
    chop_full[12][13] = 16'b00000_000000_00000;
    chop_full[12][14] = 16'b11111_111110_11111;
    chop_full[13][0] = 16'b11111_111110_11111;
    chop_full[13][1] = 16'b00000_000000_00000;
    chop_full[13][2] = 16'b00000_000000_00000;
    chop_full[13][3] = 16'b00000_000000_00000;
    chop_full[13][4] = 16'b00000_000000_00000;
    chop_full[13][5] = 16'b00000_000000_00000;
    chop_full[13][6] = 16'b00000_000000_00000;
    chop_full[13][7] = 16'b00000_000000_00000;
    chop_full[13][8] = 16'b00000_000000_00000;
    chop_full[13][9] = 16'b00000_000000_00000;
    chop_full[13][10] = 16'b00000_000000_00000;
    chop_full[13][11] = 16'b00000_000000_00000;
    chop_full[13][12] = 16'b00000_000000_00000;
    chop_full[13][13] = 16'b00000_000000_00000;
    chop_full[13][14] = 16'b11111_111110_11111;
    chop_full[14][0] = 16'b11111_111110_11111;
    chop_full[14][1] = 16'b11111_111110_11111;
    chop_full[14][2] = 16'b11111_111110_11111;
    chop_full[14][3] = 16'b11111_111110_11111;
    chop_full[14][4] = 16'b11111_111110_11111;
    chop_full[14][5] = 16'b11111_111110_11111;
    chop_full[14][6] = 16'b11111_111110_11111;
    chop_full[14][7] = 16'b11111_111110_11111;
    chop_full[14][8] = 16'b11111_111110_11111;
    chop_full[14][9] = 16'b11111_111110_11111;
    chop_full[14][10] = 16'b11111_111110_11111;
    chop_full[14][11] = 16'b11111_111110_11111;
    chop_full[14][12] = 16'b11111_111110_11111;
    chop_full[14][13] = 16'b11111_111110_11111;
    chop_full[14][14] = 16'b11111_111110_11111;
    
    end
    
    always @(posedge clk) begin
    
        prev_slow_clock <= slow_clock;
    
        case (state)
            IDLE: begin
                if (chop_ready) begin
                    state <= ANIM1;
                end
            end
            ANIM1: if (frame_tick) state <= ANIM2;
            ANIM2: if (frame_tick) state <= ANIM3;
            ANIM3: if (frame_tick) state <= ANIM4;
            ANIM4: if (frame_tick) state <= ANIM5;
            ANIM5: if (frame_tick) state <= ANIM6;
            ANIM6: if (frame_tick) state <= ANIM7;
            ANIM7: if (frame_tick) state <= ANIM8;
            ANIM8: if (frame_tick) state <= ANIM9;
            ANIM9: if (frame_tick) state <= FULL;
            FULL: begin
                //chop_ready <= 0;
                if (reset) begin
                    state <= IDLE;
                end
            end
        endcase
               
    end
    
    always @(*) begin
    
        x_idx = x - CHOPPER_TOP_LEFT_X;
        y_idx = y - CHOPPER_TOP_LEFT_Y;
        
        if (x_idx >= 0 && x_idx < 15 && y_idx >= 0 && y_idx < 15) begin
            case (state)
                IDLE: oled_data = chop_empty[y_idx][x_idx];
                ANIM1: oled_data = timing1[y_idx][x_idx];
                ANIM2: oled_data = timing2[y_idx][x_idx];
                ANIM3: oled_data = timing3[y_idx][x_idx];
                ANIM4: oled_data = timing4[y_idx][x_idx];
                ANIM5: oled_data = timing5[y_idx][x_idx];
                ANIM6: oled_data = timing6[y_idx][x_idx];
                ANIM7: oled_data = timing7[y_idx][x_idx];
                ANIM8: oled_data = timing8[y_idx][x_idx];
                ANIM9: oled_data = timing9[y_idx][x_idx];
                FULL: oled_data = chop_full[y_idx][x_idx];
                default: oled_data = chop_empty[y_idx][x_idx];
            endcase
        end else begin
            oled_data = 0;
        end
    end
    
endmodule

