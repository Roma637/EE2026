`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12.04.2025 14:24:31
// Design Name: 
// Module Name: ending_screen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ending_screen(
    input basys_clk,
    input [12:0] pixel_index,
    output reg [15:0] oled_data
);

wire [6:0] x;
wire [6:0] y;
convertToCoords coords0 (pixel_index, x, y);

reg [15:0] end_screen [0:63] [0:95] ;

initial begin
end_screen[0][0] = 16'b10001_101010_11100;
end_screen[0][1] = 16'b10001_101010_11100;
end_screen[0][2] = 16'b10001_101010_11100;
end_screen[0][3] = 16'b10001_101010_11100;
end_screen[0][4] = 16'b10001_101010_11100;
end_screen[0][5] = 16'b10001_101010_11100;
end_screen[0][6] = 16'b10001_101010_11100;
end_screen[0][7] = 16'b10001_101010_11100;
end_screen[0][8] = 16'b10001_101010_11100;
end_screen[0][9] = 16'b10001_101010_11100;
end_screen[0][10] = 16'b10001_101010_11100;
end_screen[0][11] = 16'b10001_101010_11100;
end_screen[0][12] = 16'b10001_101010_11100;
end_screen[0][13] = 16'b10001_101010_11100;
end_screen[0][14] = 16'b10001_101010_11100;
end_screen[0][15] = 16'b10001_101010_11100;
end_screen[0][16] = 16'b10001_101010_11100;
end_screen[0][17] = 16'b10001_101010_11100;
end_screen[0][18] = 16'b10001_101010_11100;
end_screen[0][19] = 16'b10001_101010_11100;
end_screen[0][20] = 16'b10001_101010_11100;
end_screen[0][21] = 16'b10001_101010_11100;
end_screen[0][22] = 16'b10001_101010_11100;
end_screen[0][23] = 16'b10001_101010_11100;
end_screen[0][24] = 16'b10001_101010_11100;
end_screen[0][25] = 16'b10001_101010_11100;
end_screen[0][26] = 16'b10001_101010_11100;
end_screen[0][27] = 16'b10001_101010_11100;
end_screen[0][28] = 16'b10001_101010_11100;
end_screen[0][29] = 16'b10001_101010_11100;
end_screen[0][30] = 16'b10001_101010_11100;
end_screen[0][31] = 16'b10001_101010_11100;
end_screen[0][32] = 16'b10001_101010_11100;
end_screen[0][33] = 16'b10001_101010_11100;
end_screen[0][34] = 16'b10001_101010_11100;
end_screen[0][35] = 16'b10001_101010_11100;
end_screen[0][36] = 16'b10001_101010_11100;
end_screen[0][37] = 16'b10001_101010_11100;
end_screen[0][38] = 16'b10001_101010_11100;
end_screen[0][39] = 16'b10001_101010_11100;
end_screen[0][40] = 16'b10001_101010_11100;
end_screen[0][41] = 16'b10001_101010_11100;
end_screen[0][42] = 16'b10001_101010_11100;
end_screen[0][43] = 16'b10001_101010_11100;
end_screen[0][44] = 16'b10001_101010_11100;
end_screen[0][45] = 16'b10001_101010_11100;
end_screen[0][46] = 16'b10001_101010_11100;
end_screen[0][47] = 16'b10001_101010_11100;
end_screen[0][48] = 16'b10001_101010_11100;
end_screen[0][49] = 16'b10001_101010_11100;
end_screen[0][50] = 16'b10001_101010_11100;
end_screen[0][51] = 16'b10001_101010_11100;
end_screen[0][52] = 16'b10001_101010_11100;
end_screen[0][53] = 16'b10001_101010_11100;
end_screen[0][54] = 16'b10001_101010_11100;
end_screen[0][55] = 16'b10001_101010_11100;
end_screen[0][56] = 16'b10001_101010_11100;
end_screen[0][57] = 16'b10001_101010_11100;
end_screen[0][58] = 16'b10001_101010_11100;
end_screen[0][59] = 16'b10001_101010_11100;
end_screen[0][60] = 16'b10001_101010_11100;
end_screen[0][61] = 16'b10001_101010_11100;
end_screen[0][62] = 16'b10001_101010_11100;
end_screen[0][63] = 16'b10001_101010_11100;
end_screen[0][64] = 16'b10001_101010_11100;
end_screen[0][65] = 16'b10001_101010_11100;
end_screen[0][66] = 16'b10001_101010_11100;
end_screen[0][67] = 16'b10001_101010_11100;
end_screen[0][68] = 16'b10001_101010_11100;
end_screen[0][69] = 16'b10001_101010_11100;
end_screen[0][70] = 16'b10001_101010_11100;
end_screen[0][71] = 16'b10001_101010_11100;
end_screen[0][72] = 16'b10001_101010_11100;
end_screen[0][73] = 16'b10001_101010_11100;
end_screen[0][74] = 16'b10001_101010_11100;
end_screen[0][75] = 16'b10001_101010_11100;
end_screen[0][76] = 16'b10001_101010_11100;
end_screen[0][77] = 16'b10001_101010_11100;
end_screen[0][78] = 16'b10001_101010_11100;
end_screen[0][79] = 16'b10001_101010_11100;
end_screen[0][80] = 16'b10001_101010_11100;
end_screen[0][81] = 16'b10001_101010_11100;
end_screen[0][82] = 16'b10001_101010_11100;
end_screen[0][83] = 16'b10001_101010_11100;
end_screen[0][84] = 16'b10001_101010_11100;
end_screen[0][85] = 16'b10001_101010_11100;
end_screen[0][86] = 16'b10001_101010_11100;
end_screen[0][87] = 16'b10001_101010_11100;
end_screen[0][88] = 16'b10001_101010_11100;
end_screen[0][89] = 16'b10001_101010_11100;
end_screen[0][90] = 16'b10001_101010_11100;
end_screen[0][91] = 16'b10001_101010_11100;
end_screen[0][92] = 16'b10001_101010_11100;
end_screen[0][93] = 16'b10001_101010_11100;
end_screen[0][94] = 16'b10001_101010_11100;
end_screen[0][95] = 16'b10001_101010_11100;
end_screen[1][0] = 16'b10001_101010_11100;
end_screen[1][1] = 16'b10001_101010_11100;
end_screen[1][2] = 16'b10001_101010_11100;
end_screen[1][3] = 16'b10001_101010_11100;
end_screen[1][4] = 16'b10001_101010_11100;
end_screen[1][5] = 16'b10001_101010_11100;
end_screen[1][6] = 16'b10001_101010_11100;
end_screen[1][7] = 16'b10001_101010_11100;
end_screen[1][8] = 16'b10001_101010_11100;
end_screen[1][9] = 16'b10001_101010_11100;
end_screen[1][10] = 16'b10001_101010_11100;
end_screen[1][11] = 16'b10001_101010_11100;
end_screen[1][12] = 16'b10001_101010_11100;
end_screen[1][13] = 16'b10001_101010_11100;
end_screen[1][14] = 16'b10001_101010_11100;
end_screen[1][15] = 16'b10001_101010_11100;
end_screen[1][16] = 16'b10001_101010_11100;
end_screen[1][17] = 16'b10001_101010_11100;
end_screen[1][18] = 16'b10001_101010_11100;
end_screen[1][19] = 16'b10001_101010_11100;
end_screen[1][20] = 16'b10001_101010_11100;
end_screen[1][21] = 16'b10001_101010_11100;
end_screen[1][22] = 16'b10001_101010_11100;
end_screen[1][23] = 16'b10001_101010_11100;
end_screen[1][24] = 16'b10001_101010_11100;
end_screen[1][25] = 16'b10001_101010_11100;
end_screen[1][26] = 16'b10001_101010_11100;
end_screen[1][27] = 16'b10001_101010_11100;
end_screen[1][28] = 16'b10001_101010_11100;
end_screen[1][29] = 16'b10001_101010_11100;
end_screen[1][30] = 16'b10001_101010_11100;
end_screen[1][31] = 16'b10001_101010_11100;
end_screen[1][32] = 16'b10001_101010_11100;
end_screen[1][33] = 16'b10001_101010_11100;
end_screen[1][34] = 16'b10001_101010_11100;
end_screen[1][35] = 16'b10001_101010_11100;
end_screen[1][36] = 16'b10001_101010_11100;
end_screen[1][37] = 16'b10001_101010_11100;
end_screen[1][38] = 16'b10001_101010_11100;
end_screen[1][39] = 16'b10001_101010_11100;
end_screen[1][40] = 16'b10001_101010_11100;
end_screen[1][41] = 16'b10001_101010_11100;
end_screen[1][42] = 16'b10001_101010_11100;
end_screen[1][43] = 16'b10001_101010_11100;
end_screen[1][44] = 16'b10001_101010_11100;
end_screen[1][45] = 16'b10001_101010_11100;
end_screen[1][46] = 16'b10001_101010_11100;
end_screen[1][47] = 16'b10001_101010_11100;
end_screen[1][48] = 16'b10001_101010_11100;
end_screen[1][49] = 16'b10001_101010_11100;
end_screen[1][50] = 16'b10001_101010_11100;
end_screen[1][51] = 16'b10001_101010_11100;
end_screen[1][52] = 16'b10001_101010_11100;
end_screen[1][53] = 16'b10001_101010_11100;
end_screen[1][54] = 16'b10001_101010_11100;
end_screen[1][55] = 16'b10001_101010_11100;
end_screen[1][56] = 16'b10001_101010_11100;
end_screen[1][57] = 16'b10001_101010_11100;
end_screen[1][58] = 16'b10001_101010_11100;
end_screen[1][59] = 16'b10001_101010_11100;
end_screen[1][60] = 16'b10001_101010_11100;
end_screen[1][61] = 16'b10001_101010_11100;
end_screen[1][62] = 16'b10001_101010_11100;
end_screen[1][63] = 16'b10001_101010_11100;
end_screen[1][64] = 16'b10001_101010_11100;
end_screen[1][65] = 16'b10001_101010_11100;
end_screen[1][66] = 16'b10001_101010_11100;
end_screen[1][67] = 16'b10001_101010_11100;
end_screen[1][68] = 16'b10001_101010_11100;
end_screen[1][69] = 16'b10001_101010_11100;
end_screen[1][70] = 16'b10001_101010_11100;
end_screen[1][71] = 16'b10001_101010_11100;
end_screen[1][72] = 16'b10001_101010_11100;
end_screen[1][73] = 16'b10001_101010_11100;
end_screen[1][74] = 16'b10001_101010_11100;
end_screen[1][75] = 16'b10001_101010_11100;
end_screen[1][76] = 16'b10001_101010_11100;
end_screen[1][77] = 16'b10001_101010_11100;
end_screen[1][78] = 16'b10001_101010_11100;
end_screen[1][79] = 16'b10001_101010_11100;
end_screen[1][80] = 16'b10001_101010_11100;
end_screen[1][81] = 16'b10001_101010_11100;
end_screen[1][82] = 16'b10001_101010_11100;
end_screen[1][83] = 16'b10001_101010_11100;
end_screen[1][84] = 16'b10001_101010_11100;
end_screen[1][85] = 16'b10001_101010_11100;
end_screen[1][86] = 16'b10001_101010_11100;
end_screen[1][87] = 16'b10001_101010_11100;
end_screen[1][88] = 16'b10001_101010_11100;
end_screen[1][89] = 16'b10001_101010_11100;
end_screen[1][90] = 16'b10001_101010_11100;
end_screen[1][91] = 16'b10001_101010_11100;
end_screen[1][92] = 16'b10001_101010_11100;
end_screen[1][93] = 16'b10001_101010_11100;
end_screen[1][94] = 16'b10001_101010_11100;
end_screen[1][95] = 16'b10001_101010_11100;
end_screen[2][0] = 16'b10001_101010_11100;
end_screen[2][1] = 16'b10001_101010_11100;
end_screen[2][2] = 16'b10001_101010_11100;
end_screen[2][3] = 16'b10001_101010_11100;
end_screen[2][4] = 16'b10001_101010_11100;
end_screen[2][5] = 16'b10001_101010_11100;
end_screen[2][6] = 16'b10001_101010_11100;
end_screen[2][7] = 16'b10001_101010_11100;
end_screen[2][8] = 16'b10001_101010_11100;
end_screen[2][9] = 16'b10001_101010_11100;
end_screen[2][10] = 16'b10001_101010_11100;
end_screen[2][11] = 16'b10001_101010_11100;
end_screen[2][12] = 16'b10001_101010_11100;
end_screen[2][13] = 16'b10001_101010_11100;
end_screen[2][14] = 16'b10001_101010_11100;
end_screen[2][15] = 16'b10001_101010_11100;
end_screen[2][16] = 16'b10001_101010_11100;
end_screen[2][17] = 16'b10001_101010_11100;
end_screen[2][18] = 16'b10001_101010_11100;
end_screen[2][19] = 16'b10001_101010_11100;
end_screen[2][20] = 16'b10001_101010_11100;
end_screen[2][21] = 16'b10001_101010_11100;
end_screen[2][22] = 16'b10001_101010_11100;
end_screen[2][23] = 16'b10001_101010_11100;
end_screen[2][24] = 16'b10001_101010_11100;
end_screen[2][25] = 16'b10001_101010_11100;
end_screen[2][26] = 16'b10001_101010_11100;
end_screen[2][27] = 16'b10001_101010_11100;
end_screen[2][28] = 16'b10001_101010_11100;
end_screen[2][29] = 16'b10001_101010_11100;
end_screen[2][30] = 16'b10001_101010_11100;
end_screen[2][31] = 16'b10001_101010_11100;
end_screen[2][32] = 16'b10001_101010_11100;
end_screen[2][33] = 16'b10001_101010_11100;
end_screen[2][34] = 16'b10001_101010_11100;
end_screen[2][35] = 16'b10001_101010_11100;
end_screen[2][36] = 16'b10001_101010_11100;
end_screen[2][37] = 16'b10001_101010_11100;
end_screen[2][38] = 16'b10001_101010_11100;
end_screen[2][39] = 16'b10001_101010_11100;
end_screen[2][40] = 16'b10001_101010_11100;
end_screen[2][41] = 16'b10001_101010_11100;
end_screen[2][42] = 16'b10001_101010_11100;
end_screen[2][43] = 16'b10001_101010_11100;
end_screen[2][44] = 16'b10001_101010_11100;
end_screen[2][45] = 16'b10001_101010_11100;
end_screen[2][46] = 16'b10001_101010_11100;
end_screen[2][47] = 16'b10001_101010_11100;
end_screen[2][48] = 16'b10001_101010_11100;
end_screen[2][49] = 16'b10001_101010_11100;
end_screen[2][50] = 16'b10001_101010_11100;
end_screen[2][51] = 16'b10001_101010_11100;
end_screen[2][52] = 16'b10001_101010_11100;
end_screen[2][53] = 16'b10001_101010_11100;
end_screen[2][54] = 16'b10001_101010_11100;
end_screen[2][55] = 16'b10001_101010_11100;
end_screen[2][56] = 16'b10001_101010_11100;
end_screen[2][57] = 16'b10001_101010_11100;
end_screen[2][58] = 16'b10001_101010_11100;
end_screen[2][59] = 16'b10001_101010_11100;
end_screen[2][60] = 16'b10001_101010_11100;
end_screen[2][61] = 16'b10001_101010_11100;
end_screen[2][62] = 16'b10001_101010_11100;
end_screen[2][63] = 16'b10001_101010_11100;
end_screen[2][64] = 16'b10001_101010_11100;
end_screen[2][65] = 16'b10001_101010_11100;
end_screen[2][66] = 16'b10001_101010_11100;
end_screen[2][67] = 16'b10001_101010_11100;
end_screen[2][68] = 16'b10001_101010_11100;
end_screen[2][69] = 16'b10001_101010_11100;
end_screen[2][70] = 16'b10001_101010_11100;
end_screen[2][71] = 16'b10001_101010_11100;
end_screen[2][72] = 16'b10001_101010_11100;
end_screen[2][73] = 16'b10001_101010_11100;
end_screen[2][74] = 16'b10001_101010_11100;
end_screen[2][75] = 16'b10001_101010_11100;
end_screen[2][76] = 16'b10001_101010_11100;
end_screen[2][77] = 16'b10001_101010_11100;
end_screen[2][78] = 16'b10001_101010_11100;
end_screen[2][79] = 16'b10001_101010_11100;
end_screen[2][80] = 16'b10001_101010_11100;
end_screen[2][81] = 16'b10001_101010_11100;
end_screen[2][82] = 16'b10001_101010_11100;
end_screen[2][83] = 16'b10001_101010_11100;
end_screen[2][84] = 16'b10001_101010_11100;
end_screen[2][85] = 16'b10001_101010_11100;
end_screen[2][86] = 16'b10001_101010_11100;
end_screen[2][87] = 16'b10001_101010_11100;
end_screen[2][88] = 16'b10001_101010_11100;
end_screen[2][89] = 16'b10001_101010_11100;
end_screen[2][90] = 16'b10001_101010_11100;
end_screen[2][91] = 16'b10001_101010_11100;
end_screen[2][92] = 16'b10001_101010_11100;
end_screen[2][93] = 16'b10001_101010_11100;
end_screen[2][94] = 16'b10001_101010_11100;
end_screen[2][95] = 16'b10001_101010_11100;
end_screen[3][0] = 16'b10001_101010_11100;
end_screen[3][1] = 16'b10001_101010_11100;
end_screen[3][2] = 16'b10001_101010_11100;
end_screen[3][3] = 16'b10001_101010_11100;
end_screen[3][4] = 16'b10001_101010_11100;
end_screen[3][5] = 16'b10001_101010_11100;
end_screen[3][6] = 16'b10001_101010_11100;
end_screen[3][7] = 16'b10001_101010_11100;
end_screen[3][8] = 16'b10001_101010_11100;
end_screen[3][9] = 16'b10001_101010_11100;
end_screen[3][10] = 16'b10001_101010_11100;
end_screen[3][11] = 16'b10001_101010_11100;
end_screen[3][12] = 16'b10001_101010_11100;
end_screen[3][13] = 16'b10001_101010_11100;
end_screen[3][14] = 16'b10001_101010_11100;
end_screen[3][15] = 16'b10001_101010_11100;
end_screen[3][16] = 16'b10001_101010_11100;
end_screen[3][17] = 16'b10001_101010_11100;
end_screen[3][18] = 16'b10001_101010_11100;
end_screen[3][19] = 16'b10001_101010_11100;
end_screen[3][20] = 16'b10001_101010_11100;
end_screen[3][21] = 16'b10001_101010_11100;
end_screen[3][22] = 16'b10001_101010_11100;
end_screen[3][23] = 16'b10001_101010_11100;
end_screen[3][24] = 16'b10001_101010_11100;
end_screen[3][25] = 16'b10001_101010_11100;
end_screen[3][26] = 16'b10001_101010_11100;
end_screen[3][27] = 16'b10001_101010_11100;
end_screen[3][28] = 16'b10001_101010_11100;
end_screen[3][29] = 16'b10000_101000_11011;
end_screen[3][30] = 16'b01000_010100_01101;
end_screen[3][31] = 16'b00100_001000_00100;
end_screen[3][32] = 16'b01000_010100_01101;
end_screen[3][33] = 16'b10001_101010_11100;
end_screen[3][34] = 16'b10001_101010_11100;
end_screen[3][35] = 16'b10001_101010_11100;
end_screen[3][36] = 16'b10001_101010_11100;
end_screen[3][37] = 16'b10001_101010_11100;
end_screen[3][38] = 16'b10001_101010_11100;
end_screen[3][39] = 16'b10001_101010_11100;
end_screen[3][40] = 16'b10001_101010_11100;
end_screen[3][41] = 16'b10001_101010_11100;
end_screen[3][42] = 16'b10001_101010_11100;
end_screen[3][43] = 16'b10001_101010_11100;
end_screen[3][44] = 16'b10001_101010_11100;
end_screen[3][45] = 16'b10001_101010_11100;
end_screen[3][46] = 16'b10001_101010_11100;
end_screen[3][47] = 16'b10001_101010_11100;
end_screen[3][48] = 16'b10001_101010_11100;
end_screen[3][49] = 16'b01111_100101_11001;
end_screen[3][50] = 16'b00110_001111_01001;
end_screen[3][51] = 16'b00100_001000_00100;
end_screen[3][52] = 16'b01100_011101_10011;
end_screen[3][53] = 16'b10001_101010_11100;
end_screen[3][54] = 16'b10001_101010_11100;
end_screen[3][55] = 16'b10001_101010_11100;
end_screen[3][56] = 16'b10001_101010_11100;
end_screen[3][57] = 16'b10001_101010_11100;
end_screen[3][58] = 16'b10001_101010_11100;
end_screen[3][59] = 16'b10001_101010_11100;
end_screen[3][60] = 16'b10001_101010_11100;
end_screen[3][61] = 16'b10001_101010_11100;
end_screen[3][62] = 16'b10001_101010_11100;
end_screen[3][63] = 16'b10001_101010_11100;
end_screen[3][64] = 16'b10001_101010_11100;
end_screen[3][65] = 16'b10001_101010_11100;
end_screen[3][66] = 16'b10001_101010_11100;
end_screen[3][67] = 16'b10001_101010_11100;
end_screen[3][68] = 16'b10001_101010_11100;
end_screen[3][69] = 16'b10001_101010_11100;
end_screen[3][70] = 16'b10001_101010_11100;
end_screen[3][71] = 16'b10001_101010_11100;
end_screen[3][72] = 16'b10001_101010_11100;
end_screen[3][73] = 16'b10001_101010_11100;
end_screen[3][74] = 16'b10001_101010_11100;
end_screen[3][75] = 16'b10001_101010_11100;
end_screen[3][76] = 16'b10001_101010_11100;
end_screen[3][77] = 16'b10001_101010_11100;
end_screen[3][78] = 16'b10001_101010_11100;
end_screen[3][79] = 16'b10001_101010_11100;
end_screen[3][80] = 16'b10001_101010_11100;
end_screen[3][81] = 16'b10001_101010_11100;
end_screen[3][82] = 16'b10001_101010_11100;
end_screen[3][83] = 16'b10001_101010_11100;
end_screen[3][84] = 16'b10001_101010_11100;
end_screen[3][85] = 16'b10001_101010_11100;
end_screen[3][86] = 16'b10001_101010_11100;
end_screen[3][87] = 16'b10001_101010_11100;
end_screen[3][88] = 16'b10001_101010_11100;
end_screen[3][89] = 16'b10001_101010_11100;
end_screen[3][90] = 16'b10001_101010_11100;
end_screen[3][91] = 16'b10001_101010_11100;
end_screen[3][92] = 16'b10001_101010_11100;
end_screen[3][93] = 16'b10001_101010_11100;
end_screen[3][94] = 16'b10001_101010_11100;
end_screen[3][95] = 16'b10001_101010_11100;
end_screen[4][0] = 16'b10001_101010_11100;
end_screen[4][1] = 16'b10001_101010_11100;
end_screen[4][2] = 16'b10001_101010_11100;
end_screen[4][3] = 16'b10001_101010_11100;
end_screen[4][4] = 16'b10001_101010_11100;
end_screen[4][5] = 16'b10001_101010_11100;
end_screen[4][6] = 16'b10001_101010_11100;
end_screen[4][7] = 16'b10001_101010_11100;
end_screen[4][8] = 16'b10001_101010_11100;
end_screen[4][9] = 16'b10001_101010_11100;
end_screen[4][10] = 16'b10001_101010_11100;
end_screen[4][11] = 16'b10001_101010_11100;
end_screen[4][12] = 16'b10001_101010_11100;
end_screen[4][13] = 16'b10001_101010_11100;
end_screen[4][14] = 16'b10001_101010_11100;
end_screen[4][15] = 16'b10001_101010_11100;
end_screen[4][16] = 16'b10001_101010_11100;
end_screen[4][17] = 16'b10001_101010_11100;
end_screen[4][18] = 16'b10001_101010_11100;
end_screen[4][19] = 16'b10001_101010_11100;
end_screen[4][20] = 16'b10001_101010_11100;
end_screen[4][21] = 16'b10001_101010_11100;
end_screen[4][22] = 16'b10001_101010_11100;
end_screen[4][23] = 16'b10001_101010_11100;
end_screen[4][24] = 16'b10001_101010_11100;
end_screen[4][25] = 16'b10001_101010_11100;
end_screen[4][26] = 16'b10001_101010_11100;
end_screen[4][27] = 16'b10001_101010_11100;
end_screen[4][28] = 16'b10001_101010_11100;
end_screen[4][29] = 16'b01011_011011_10010;
end_screen[4][30] = 16'b00100_001000_00100;
end_screen[4][31] = 16'b00100_001000_00100;
end_screen[4][32] = 16'b00100_001000_00100;
end_screen[4][33] = 16'b01100_011101_10011;
end_screen[4][34] = 16'b10001_101010_11100;
end_screen[4][35] = 16'b10001_101010_11100;
end_screen[4][36] = 16'b10001_101010_11100;
end_screen[4][37] = 16'b10001_101010_11100;
end_screen[4][38] = 16'b10001_101010_11100;
end_screen[4][39] = 16'b10001_101010_11100;
end_screen[4][40] = 16'b10001_101010_11100;
end_screen[4][41] = 16'b10001_101010_11100;
end_screen[4][42] = 16'b10001_101010_11100;
end_screen[4][43] = 16'b10001_101010_11100;
end_screen[4][44] = 16'b10001_101010_11100;
end_screen[4][45] = 16'b10001_101010_11100;
end_screen[4][46] = 16'b10001_101010_11100;
end_screen[4][47] = 16'b10001_101010_11100;
end_screen[4][48] = 16'b10001_101010_11100;
end_screen[4][49] = 16'b00111_010001_01011;
end_screen[4][50] = 16'b00100_001000_00100;
end_screen[4][51] = 16'b00100_001000_00100;
end_screen[4][52] = 16'b00100_001000_00100;
end_screen[4][53] = 16'b01110_100011_10111;
end_screen[4][54] = 16'b10001_101010_11100;
end_screen[4][55] = 16'b10001_101010_11100;
end_screen[4][56] = 16'b10001_101010_11100;
end_screen[4][57] = 16'b10001_101010_11100;
end_screen[4][58] = 16'b10001_101010_11100;
end_screen[4][59] = 16'b10001_101010_11100;
end_screen[4][60] = 16'b10001_101010_11100;
end_screen[4][61] = 16'b10001_101010_11100;
end_screen[4][62] = 16'b10001_101010_11100;
end_screen[4][63] = 16'b10001_101010_11100;
end_screen[4][64] = 16'b10001_101010_11100;
end_screen[4][65] = 16'b10001_101010_11100;
end_screen[4][66] = 16'b10001_101010_11100;
end_screen[4][67] = 16'b01110_100011_10111;
end_screen[4][68] = 16'b00101_001011_00111;
end_screen[4][69] = 16'b00100_001000_00100;
end_screen[4][70] = 16'b01100_011101_10011;
end_screen[4][71] = 16'b10001_101010_11100;
end_screen[4][72] = 16'b10001_101010_11100;
end_screen[4][73] = 16'b10001_101010_11100;
end_screen[4][74] = 16'b10001_101010_11100;
end_screen[4][75] = 16'b10001_101010_11100;
end_screen[4][76] = 16'b10001_101010_11100;
end_screen[4][77] = 16'b10001_101010_11100;
end_screen[4][78] = 16'b10001_101010_11100;
end_screen[4][79] = 16'b10001_101010_11100;
end_screen[4][80] = 16'b10001_101010_11100;
end_screen[4][81] = 16'b10001_101010_11100;
end_screen[4][82] = 16'b10001_101010_11100;
end_screen[4][83] = 16'b10001_101010_11100;
end_screen[4][84] = 16'b10001_101010_11100;
end_screen[4][85] = 16'b10001_101010_11100;
end_screen[4][86] = 16'b10001_101010_11100;
end_screen[4][87] = 16'b10001_101010_11100;
end_screen[4][88] = 16'b10001_101010_11100;
end_screen[4][89] = 16'b10001_101010_11100;
end_screen[4][90] = 16'b10001_101010_11100;
end_screen[4][91] = 16'b10001_101010_11100;
end_screen[4][92] = 16'b10001_101010_11100;
end_screen[4][93] = 16'b10001_101010_11100;
end_screen[4][94] = 16'b10001_101010_11100;
end_screen[4][95] = 16'b10001_101010_11100;
end_screen[5][0] = 16'b10001_101010_11100;
end_screen[5][1] = 16'b10001_101010_11100;
end_screen[5][2] = 16'b10001_101010_11100;
end_screen[5][3] = 16'b10001_101010_11100;
end_screen[5][4] = 16'b10001_101010_11100;
end_screen[5][5] = 16'b10001_101010_11100;
end_screen[5][6] = 16'b10001_101010_11100;
end_screen[5][7] = 16'b10001_101010_11100;
end_screen[5][8] = 16'b10001_101010_11100;
end_screen[5][9] = 16'b10001_101010_11100;
end_screen[5][10] = 16'b10001_101010_11100;
end_screen[5][11] = 16'b10001_101010_11100;
end_screen[5][12] = 16'b10001_101010_11100;
end_screen[5][13] = 16'b10001_101010_11100;
end_screen[5][14] = 16'b10001_101010_11100;
end_screen[5][15] = 16'b10001_101010_11100;
end_screen[5][16] = 16'b10001_101010_11100;
end_screen[5][17] = 16'b10001_101010_11100;
end_screen[5][18] = 16'b10000_101000_11011;
end_screen[5][19] = 16'b01000_010100_01101;
end_screen[5][20] = 16'b00100_001000_00100;
end_screen[5][21] = 16'b00100_001000_00100;
end_screen[5][22] = 16'b00100_001000_00100;
end_screen[5][23] = 16'b00100_001000_00100;
end_screen[5][24] = 16'b00100_001000_00100;
end_screen[5][25] = 16'b00100_001000_00100;
end_screen[5][26] = 16'b00111_010001_01011;
end_screen[5][27] = 16'b10000_100111_11010;
end_screen[5][28] = 16'b10001_101010_11100;
end_screen[5][29] = 16'b01000_010100_01101;
end_screen[5][30] = 16'b00100_001000_00100;
end_screen[5][31] = 16'b00100_001000_00100;
end_screen[5][32] = 16'b00100_001000_00100;
end_screen[5][33] = 16'b01000_010100_01101;
end_screen[5][34] = 16'b10001_101010_11100;
end_screen[5][35] = 16'b10001_101010_11100;
end_screen[5][36] = 16'b10001_101010_11100;
end_screen[5][37] = 16'b10001_101010_11100;
end_screen[5][38] = 16'b10001_101010_11100;
end_screen[5][39] = 16'b10001_101010_11100;
end_screen[5][40] = 16'b10001_101010_11100;
end_screen[5][41] = 16'b10001_101010_11100;
end_screen[5][42] = 16'b10001_101010_11100;
end_screen[5][43] = 16'b10001_101010_11100;
end_screen[5][44] = 16'b10001_101010_11100;
end_screen[5][45] = 16'b10001_101010_11100;
end_screen[5][46] = 16'b10001_101010_11100;
end_screen[5][47] = 16'b10001_101010_11100;
end_screen[5][48] = 16'b10001_101010_11100;
end_screen[5][49] = 16'b00100_001000_00100;
end_screen[5][50] = 16'b00100_001000_00100;
end_screen[5][51] = 16'b00100_001000_00100;
end_screen[5][52] = 16'b00100_001000_00100;
end_screen[5][53] = 16'b01100_011101_10011;
end_screen[5][54] = 16'b10001_101010_11100;
end_screen[5][55] = 16'b10001_101010_11100;
end_screen[5][56] = 16'b10001_101010_11100;
end_screen[5][57] = 16'b10001_101010_11100;
end_screen[5][58] = 16'b10001_101010_11100;
end_screen[5][59] = 16'b10001_101010_11100;
end_screen[5][60] = 16'b10001_101010_11100;
end_screen[5][61] = 16'b10001_101010_11100;
end_screen[5][62] = 16'b10001_101010_11100;
end_screen[5][63] = 16'b10001_101010_11100;
end_screen[5][64] = 16'b10001_101010_11100;
end_screen[5][65] = 16'b10001_101010_11100;
end_screen[5][66] = 16'b10001_101010_11100;
end_screen[5][67] = 16'b00110_001111_01001;
end_screen[5][68] = 16'b00100_001000_00100;
end_screen[5][69] = 16'b00100_001000_00100;
end_screen[5][70] = 16'b00100_001000_00100;
end_screen[5][71] = 16'b01111_100101_11001;
end_screen[5][72] = 16'b10001_101010_11100;
end_screen[5][73] = 16'b10001_101010_11100;
end_screen[5][74] = 16'b10001_101010_11100;
end_screen[5][75] = 16'b10001_101010_11100;
end_screen[5][76] = 16'b10001_101010_11100;
end_screen[5][77] = 16'b10001_101010_11100;
end_screen[5][78] = 16'b10001_101010_11100;
end_screen[5][79] = 16'b10001_101010_11100;
end_screen[5][80] = 16'b10001_101010_11100;
end_screen[5][81] = 16'b10001_101010_11100;
end_screen[5][82] = 16'b10001_101010_11100;
end_screen[5][83] = 16'b10001_101010_11100;
end_screen[5][84] = 16'b10001_101010_11100;
end_screen[5][85] = 16'b10001_101010_11100;
end_screen[5][86] = 16'b10001_101010_11100;
end_screen[5][87] = 16'b10001_101010_11100;
end_screen[5][88] = 16'b10001_101010_11100;
end_screen[5][89] = 16'b10001_101010_11100;
end_screen[5][90] = 16'b10001_101010_11100;
end_screen[5][91] = 16'b10001_101010_11100;
end_screen[5][92] = 16'b10001_101010_11100;
end_screen[5][93] = 16'b10001_101010_11100;
end_screen[5][94] = 16'b10001_101010_11100;
end_screen[5][95] = 16'b10001_101010_11100;
end_screen[6][0] = 16'b10001_101010_11100;
end_screen[6][1] = 16'b10001_101010_11100;
end_screen[6][2] = 16'b10001_101010_11100;
end_screen[6][3] = 16'b10001_101010_11100;
end_screen[6][4] = 16'b10001_101010_11100;
end_screen[6][5] = 16'b10001_101010_11100;
end_screen[6][6] = 16'b10001_101010_11100;
end_screen[6][7] = 16'b10001_101010_11100;
end_screen[6][8] = 16'b10001_101010_11100;
end_screen[6][9] = 16'b10001_101010_11100;
end_screen[6][10] = 16'b10001_101010_11100;
end_screen[6][11] = 16'b10001_101010_11100;
end_screen[6][12] = 16'b10001_101010_11100;
end_screen[6][13] = 16'b10001_101010_11100;
end_screen[6][14] = 16'b10001_101010_11100;
end_screen[6][15] = 16'b10001_101010_11100;
end_screen[6][16] = 16'b10001_101010_11100;
end_screen[6][17] = 16'b10001_101010_11100;
end_screen[6][18] = 16'b01011_011011_10010;
end_screen[6][19] = 16'b00100_001000_00100;
end_screen[6][20] = 16'b00100_001000_00100;
end_screen[6][21] = 16'b00100_001000_00100;
end_screen[6][22] = 16'b00100_001000_00100;
end_screen[6][23] = 16'b00100_001000_00100;
end_screen[6][24] = 16'b00100_001000_00100;
end_screen[6][25] = 16'b00100_001000_00100;
end_screen[6][26] = 16'b00100_001000_00100;
end_screen[6][27] = 16'b01011_011011_10010;
end_screen[6][28] = 16'b10001_101010_11100;
end_screen[6][29] = 16'b01011_011011_10010;
end_screen[6][30] = 16'b00100_001000_00100;
end_screen[6][31] = 16'b00100_001000_00100;
end_screen[6][32] = 16'b00100_001000_00100;
end_screen[6][33] = 16'b01100_011101_10011;
end_screen[6][34] = 16'b10001_101010_11100;
end_screen[6][35] = 16'b10001_101010_11100;
end_screen[6][36] = 16'b10001_101010_11100;
end_screen[6][37] = 16'b10001_101010_11100;
end_screen[6][38] = 16'b10001_101010_11100;
end_screen[6][39] = 16'b10001_101010_11100;
end_screen[6][40] = 16'b10001_101010_11100;
end_screen[6][41] = 16'b10001_101010_11100;
end_screen[6][42] = 16'b10001_101010_11100;
end_screen[6][43] = 16'b10001_101010_11100;
end_screen[6][44] = 16'b10001_101010_11100;
end_screen[6][45] = 16'b10001_101010_11100;
end_screen[6][46] = 16'b10001_101010_11100;
end_screen[6][47] = 16'b10001_101010_11100;
end_screen[6][48] = 16'b10001_101010_11100;
end_screen[6][49] = 16'b00111_010001_01011;
end_screen[6][50] = 16'b00100_001000_00100;
end_screen[6][51] = 16'b00100_001000_00100;
end_screen[6][52] = 16'b00100_001000_00100;
end_screen[6][53] = 16'b01110_100011_10111;
end_screen[6][54] = 16'b10001_101010_11100;
end_screen[6][55] = 16'b10001_101010_11100;
end_screen[6][56] = 16'b10001_101010_11100;
end_screen[6][57] = 16'b10001_101010_11100;
end_screen[6][58] = 16'b10001_101010_11100;
end_screen[6][59] = 16'b10001_101010_11100;
end_screen[6][60] = 16'b10001_101010_11100;
end_screen[6][61] = 16'b10001_101010_11100;
end_screen[6][62] = 16'b10001_101010_11100;
end_screen[6][63] = 16'b10001_101010_11100;
end_screen[6][64] = 16'b10001_101010_11100;
end_screen[6][65] = 16'b10001_101010_11100;
end_screen[6][66] = 16'b10001_101010_11100;
end_screen[6][67] = 16'b00100_001000_00100;
end_screen[6][68] = 16'b00100_001000_00100;
end_screen[6][69] = 16'b00100_001000_00100;
end_screen[6][70] = 16'b00100_001000_00100;
end_screen[6][71] = 16'b01110_100011_10111;
end_screen[6][72] = 16'b10001_101010_11100;
end_screen[6][73] = 16'b10001_101010_11100;
end_screen[6][74] = 16'b10001_101010_11100;
end_screen[6][75] = 16'b10001_101010_11100;
end_screen[6][76] = 16'b10001_101010_11100;
end_screen[6][77] = 16'b10001_101010_11100;
end_screen[6][78] = 16'b10001_101010_11100;
end_screen[6][79] = 16'b10001_101010_11100;
end_screen[6][80] = 16'b10001_101010_11100;
end_screen[6][81] = 16'b10001_101010_11100;
end_screen[6][82] = 16'b10001_101010_11100;
end_screen[6][83] = 16'b10001_101010_11100;
end_screen[6][84] = 16'b10001_101010_11100;
end_screen[6][85] = 16'b10001_101010_11100;
end_screen[6][86] = 16'b10001_101010_11100;
end_screen[6][87] = 16'b10001_101010_11100;
end_screen[6][88] = 16'b10001_101010_11100;
end_screen[6][89] = 16'b10001_101010_11100;
end_screen[6][90] = 16'b10001_101010_11100;
end_screen[6][91] = 16'b10001_101010_11100;
end_screen[6][92] = 16'b10001_101010_11100;
end_screen[6][93] = 16'b10001_101010_11100;
end_screen[6][94] = 16'b10001_101010_11100;
end_screen[6][95] = 16'b10001_101010_11100;
end_screen[7][0] = 16'b10001_101010_11100;
end_screen[7][1] = 16'b10001_101010_11100;
end_screen[7][2] = 16'b10001_101010_11100;
end_screen[7][3] = 16'b10001_101010_11100;
end_screen[7][4] = 16'b10001_101010_11100;
end_screen[7][5] = 16'b10001_101010_11100;
end_screen[7][6] = 16'b10001_101010_11100;
end_screen[7][7] = 16'b10001_101010_11100;
end_screen[7][8] = 16'b10001_101010_11100;
end_screen[7][9] = 16'b10001_101010_11100;
end_screen[7][10] = 16'b10001_101010_11100;
end_screen[7][11] = 16'b10001_101010_11100;
end_screen[7][12] = 16'b10001_101010_11100;
end_screen[7][13] = 16'b10001_101010_11100;
end_screen[7][14] = 16'b10001_101010_11100;
end_screen[7][15] = 16'b10001_101010_11100;
end_screen[7][16] = 16'b10001_101010_11100;
end_screen[7][17] = 16'b10001_101010_11100;
end_screen[7][18] = 16'b01000_010100_01101;
end_screen[7][19] = 16'b00100_001000_00100;
end_screen[7][20] = 16'b00100_001000_00100;
end_screen[7][21] = 16'b00100_001000_00100;
end_screen[7][22] = 16'b00100_001000_00100;
end_screen[7][23] = 16'b00100_001000_00100;
end_screen[7][24] = 16'b00100_001000_00100;
end_screen[7][25] = 16'b00100_001000_00100;
end_screen[7][26] = 16'b00100_001000_00100;
end_screen[7][27] = 16'b01011_011011_10010;
end_screen[7][28] = 16'b10001_101010_11100;
end_screen[7][29] = 16'b10000_101000_11011;
end_screen[7][30] = 16'b01000_010100_01101;
end_screen[7][31] = 16'b00100_001000_00100;
end_screen[7][32] = 16'b01000_010100_01101;
end_screen[7][33] = 16'b10000_101000_11011;
end_screen[7][34] = 16'b10001_101010_11100;
end_screen[7][35] = 16'b10001_101010_11100;
end_screen[7][36] = 16'b10001_101010_11100;
end_screen[7][37] = 16'b10001_101010_11100;
end_screen[7][38] = 16'b10001_101010_11100;
end_screen[7][39] = 16'b10001_101010_11100;
end_screen[7][40] = 16'b10001_101010_11100;
end_screen[7][41] = 16'b10001_101010_11100;
end_screen[7][42] = 16'b10001_101010_11100;
end_screen[7][43] = 16'b10001_101010_11100;
end_screen[7][44] = 16'b10001_101010_11100;
end_screen[7][45] = 16'b10001_101010_11100;
end_screen[7][46] = 16'b10001_101010_11100;
end_screen[7][47] = 16'b10001_101010_11100;
end_screen[7][48] = 16'b10001_101010_11100;
end_screen[7][49] = 16'b01111_100101_11001;
end_screen[7][50] = 16'b00110_001111_01001;
end_screen[7][51] = 16'b00100_001000_00100;
end_screen[7][52] = 16'b01011_011011_10010;
end_screen[7][53] = 16'b10001_101010_11100;
end_screen[7][54] = 16'b10001_101010_11100;
end_screen[7][55] = 16'b10001_101010_11100;
end_screen[7][56] = 16'b10001_101010_11100;
end_screen[7][57] = 16'b10001_101010_11100;
end_screen[7][58] = 16'b10001_101010_11100;
end_screen[7][59] = 16'b10001_101010_11100;
end_screen[7][60] = 16'b10001_101010_11100;
end_screen[7][61] = 16'b10001_101010_11100;
end_screen[7][62] = 16'b10001_101010_11100;
end_screen[7][63] = 16'b10001_101010_11100;
end_screen[7][64] = 16'b10001_101010_11100;
end_screen[7][65] = 16'b10001_101010_11100;
end_screen[7][66] = 16'b10001_101010_11100;
end_screen[7][67] = 16'b00100_001000_00100;
end_screen[7][68] = 16'b00100_001000_00100;
end_screen[7][69] = 16'b00100_001000_00100;
end_screen[7][70] = 16'b00100_001000_00100;
end_screen[7][71] = 16'b01110_100011_10111;
end_screen[7][72] = 16'b10001_101010_11100;
end_screen[7][73] = 16'b10001_101010_11100;
end_screen[7][74] = 16'b10001_101010_11100;
end_screen[7][75] = 16'b10001_101010_11100;
end_screen[7][76] = 16'b10001_101010_11100;
end_screen[7][77] = 16'b10001_101010_11100;
end_screen[7][78] = 16'b10001_101010_11100;
end_screen[7][79] = 16'b10001_101010_11100;
end_screen[7][80] = 16'b10001_101010_11100;
end_screen[7][81] = 16'b10001_101010_11100;
end_screen[7][82] = 16'b10001_101010_11100;
end_screen[7][83] = 16'b10001_101010_11100;
end_screen[7][84] = 16'b10001_101010_11100;
end_screen[7][85] = 16'b10001_101010_11100;
end_screen[7][86] = 16'b10001_101010_11100;
end_screen[7][87] = 16'b10001_101010_11100;
end_screen[7][88] = 16'b10001_101010_11100;
end_screen[7][89] = 16'b10001_101010_11100;
end_screen[7][90] = 16'b10001_101010_11100;
end_screen[7][91] = 16'b10001_101010_11100;
end_screen[7][92] = 16'b10001_101010_11100;
end_screen[7][93] = 16'b10001_101010_11100;
end_screen[7][94] = 16'b10001_101010_11100;
end_screen[7][95] = 16'b10001_101010_11100;
end_screen[8][0] = 16'b10001_101010_11100;
end_screen[8][1] = 16'b10001_101010_11100;
end_screen[8][2] = 16'b10001_101010_11100;
end_screen[8][3] = 16'b10001_101010_11100;
end_screen[8][4] = 16'b10001_101010_11100;
end_screen[8][5] = 16'b10001_101010_11100;
end_screen[8][6] = 16'b10001_101010_11100;
end_screen[8][7] = 16'b10001_101010_11100;
end_screen[8][8] = 16'b10001_101010_11100;
end_screen[8][9] = 16'b10001_101010_11100;
end_screen[8][10] = 16'b10001_101010_11100;
end_screen[8][11] = 16'b10001_101010_11100;
end_screen[8][12] = 16'b10001_101010_11100;
end_screen[8][13] = 16'b10001_101010_11100;
end_screen[8][14] = 16'b10001_101010_11100;
end_screen[8][15] = 16'b10001_101010_11100;
end_screen[8][16] = 16'b10001_101010_11100;
end_screen[8][17] = 16'b10001_101010_11100;
end_screen[8][18] = 16'b01000_010100_01101;
end_screen[8][19] = 16'b00100_001000_00100;
end_screen[8][20] = 16'b00100_001000_00100;
end_screen[8][21] = 16'b00100_001000_00100;
end_screen[8][22] = 16'b00100_001000_00100;
end_screen[8][23] = 16'b00100_001000_00100;
end_screen[8][24] = 16'b00100_001000_00100;
end_screen[8][25] = 16'b00100_001000_00100;
end_screen[8][26] = 16'b00111_010001_01011;
end_screen[8][27] = 16'b10000_100111_11010;
end_screen[8][28] = 16'b10001_101010_11100;
end_screen[8][29] = 16'b10001_101010_11100;
end_screen[8][30] = 16'b01101_011111_10101;
end_screen[8][31] = 16'b01100_011101_10011;
end_screen[8][32] = 16'b01101_011111_10101;
end_screen[8][33] = 16'b10001_101010_11100;
end_screen[8][34] = 16'b10001_101010_11100;
end_screen[8][35] = 16'b10001_101010_11100;
end_screen[8][36] = 16'b10001_101010_11100;
end_screen[8][37] = 16'b10001_101010_11100;
end_screen[8][38] = 16'b10001_101010_11100;
end_screen[8][39] = 16'b10001_101010_11100;
end_screen[8][40] = 16'b10001_101010_11100;
end_screen[8][41] = 16'b10001_101010_11100;
end_screen[8][42] = 16'b10001_101010_11100;
end_screen[8][43] = 16'b10001_101010_11100;
end_screen[8][44] = 16'b10001_101010_11100;
end_screen[8][45] = 16'b10001_101010_11100;
end_screen[8][46] = 16'b10001_101010_11100;
end_screen[8][47] = 16'b10001_101010_11100;
end_screen[8][48] = 16'b10001_101010_11100;
end_screen[8][49] = 16'b10001_101010_11100;
end_screen[8][50] = 16'b01100_011101_10011;
end_screen[8][51] = 16'b01100_011101_10011;
end_screen[8][52] = 16'b01110_100011_10111;
end_screen[8][53] = 16'b10001_101010_11100;
end_screen[8][54] = 16'b10001_101010_11100;
end_screen[8][55] = 16'b10001_101010_11100;
end_screen[8][56] = 16'b10001_101010_11100;
end_screen[8][57] = 16'b10001_101010_11100;
end_screen[8][58] = 16'b01101_011111_10101;
end_screen[8][59] = 16'b01100_011101_10011;
end_screen[8][60] = 16'b01100_011101_10011;
end_screen[8][61] = 16'b01100_011101_10011;
end_screen[8][62] = 16'b01100_011101_10011;
end_screen[8][63] = 16'b10000_101000_11011;
end_screen[8][64] = 16'b10001_101010_11100;
end_screen[8][65] = 16'b10001_101010_11100;
end_screen[8][66] = 16'b10001_101010_11100;
end_screen[8][67] = 16'b00100_001000_00100;
end_screen[8][68] = 16'b00100_001000_00100;
end_screen[8][69] = 16'b00100_001000_00100;
end_screen[8][70] = 16'b00100_001000_00100;
end_screen[8][71] = 16'b01110_100011_10111;
end_screen[8][72] = 16'b01100_011101_10011;
end_screen[8][73] = 16'b01100_011101_10011;
end_screen[8][74] = 16'b01100_011101_10011;
end_screen[8][75] = 16'b01110_100011_10111;
end_screen[8][76] = 16'b10001_101010_11100;
end_screen[8][77] = 16'b10001_101010_11100;
end_screen[8][78] = 16'b10001_101010_11100;
end_screen[8][79] = 16'b10001_101010_11100;
end_screen[8][80] = 16'b10001_101010_11100;
end_screen[8][81] = 16'b10001_101010_11100;
end_screen[8][82] = 16'b10001_101010_11100;
end_screen[8][83] = 16'b10001_101010_11100;
end_screen[8][84] = 16'b10001_101010_11100;
end_screen[8][85] = 16'b10001_101010_11100;
end_screen[8][86] = 16'b10001_101010_11100;
end_screen[8][87] = 16'b10001_101010_11100;
end_screen[8][88] = 16'b10001_101010_11100;
end_screen[8][89] = 16'b10001_101010_11100;
end_screen[8][90] = 16'b10001_101010_11100;
end_screen[8][91] = 16'b10001_101010_11100;
end_screen[8][92] = 16'b10001_101010_11100;
end_screen[8][93] = 16'b10001_101010_11100;
end_screen[8][94] = 16'b10001_101010_11100;
end_screen[8][95] = 16'b10001_101010_11100;
end_screen[9][0] = 16'b10001_101010_11100;
end_screen[9][1] = 16'b10001_101010_11100;
end_screen[9][2] = 16'b10001_101010_11100;
end_screen[9][3] = 16'b10001_101010_11100;
end_screen[9][4] = 16'b10001_101010_11100;
end_screen[9][5] = 16'b10001_101010_11100;
end_screen[9][6] = 16'b10001_101010_11100;
end_screen[9][7] = 16'b10001_101010_11100;
end_screen[9][8] = 16'b10001_101010_11100;
end_screen[9][9] = 16'b10001_101010_11100;
end_screen[9][10] = 16'b10001_101010_11100;
end_screen[9][11] = 16'b10001_101010_11100;
end_screen[9][12] = 16'b10001_101010_11100;
end_screen[9][13] = 16'b10001_101010_11100;
end_screen[9][14] = 16'b10001_101010_11100;
end_screen[9][15] = 16'b10001_101010_11100;
end_screen[9][16] = 16'b10001_101010_11100;
end_screen[9][17] = 16'b10001_101010_11100;
end_screen[9][18] = 16'b01000_010100_01101;
end_screen[9][19] = 16'b00100_001000_00100;
end_screen[9][20] = 16'b00100_001000_00100;
end_screen[9][21] = 16'b00100_001000_00100;
end_screen[9][22] = 16'b01000_010100_01101;
end_screen[9][23] = 16'b10001_101010_11100;
end_screen[9][24] = 16'b10001_101010_11100;
end_screen[9][25] = 16'b10001_101010_11100;
end_screen[9][26] = 16'b10001_101010_11100;
end_screen[9][27] = 16'b10001_101010_11100;
end_screen[9][28] = 16'b10001_101010_11100;
end_screen[9][29] = 16'b01101_011111_10101;
end_screen[9][30] = 16'b00100_001000_00100;
end_screen[9][31] = 16'b00100_001000_00100;
end_screen[9][32] = 16'b00100_001000_00100;
end_screen[9][33] = 16'b01101_011111_10101;
end_screen[9][34] = 16'b10001_101010_11100;
end_screen[9][35] = 16'b10001_101010_11100;
end_screen[9][36] = 16'b01110_100011_10111;
end_screen[9][37] = 16'b00101_001011_00111;
end_screen[9][38] = 16'b00111_010001_01011;
end_screen[9][39] = 16'b01110_100011_10111;
end_screen[9][40] = 16'b01100_011101_10011;
end_screen[9][41] = 16'b00101_001011_00111;
end_screen[9][42] = 16'b00100_001000_00100;
end_screen[9][43] = 16'b00100_001000_00100;
end_screen[9][44] = 16'b01011_011011_10010;
end_screen[9][45] = 16'b10000_101000_11011;
end_screen[9][46] = 16'b10001_101010_11100;
end_screen[9][47] = 16'b10001_101010_11100;
end_screen[9][48] = 16'b10001_101010_11100;
end_screen[9][49] = 16'b01010_011001_10000;
end_screen[9][50] = 16'b00100_001000_00100;
end_screen[9][51] = 16'b00100_001000_00100;
end_screen[9][52] = 16'b00100_001000_00100;
end_screen[9][53] = 16'b10000_100111_11010;
end_screen[9][54] = 16'b10001_101010_11100;
end_screen[9][55] = 16'b10001_101010_11100;
end_screen[9][56] = 16'b10000_100111_11010;
end_screen[9][57] = 16'b00111_010001_01011;
end_screen[9][58] = 16'b00100_001000_00100;
end_screen[9][59] = 16'b00100_001000_00100;
end_screen[9][60] = 16'b00100_001000_00100;
end_screen[9][61] = 16'b00100_001000_00100;
end_screen[9][62] = 16'b00100_001000_00100;
end_screen[9][63] = 16'b00100_001000_00100;
end_screen[9][64] = 16'b01101_100001_10110;
end_screen[9][65] = 16'b10001_101010_11100;
end_screen[9][66] = 16'b10001_101010_11100;
end_screen[9][67] = 16'b00100_001000_00100;
end_screen[9][68] = 16'b00100_001000_00100;
end_screen[9][69] = 16'b00100_001000_00100;
end_screen[9][70] = 16'b00100_001000_00100;
end_screen[9][71] = 16'b00100_001000_00100;
end_screen[9][72] = 16'b00100_001000_00100;
end_screen[9][73] = 16'b00100_001000_00100;
end_screen[9][74] = 16'b00100_001000_00100;
end_screen[9][75] = 16'b00100_001000_00100;
end_screen[9][76] = 16'b01010_011001_10000;
end_screen[9][77] = 16'b10001_101010_11100;
end_screen[9][78] = 16'b10001_101010_11100;
end_screen[9][79] = 16'b10001_101010_11100;
end_screen[9][80] = 16'b10001_101010_11100;
end_screen[9][81] = 16'b10001_101010_11100;
end_screen[9][82] = 16'b10001_101010_11100;
end_screen[9][83] = 16'b10001_101010_11100;
end_screen[9][84] = 16'b10001_101010_11100;
end_screen[9][85] = 16'b10001_101010_11100;
end_screen[9][86] = 16'b10001_101010_11100;
end_screen[9][87] = 16'b10001_101010_11100;
end_screen[9][88] = 16'b10001_101010_11100;
end_screen[9][89] = 16'b10001_101010_11100;
end_screen[9][90] = 16'b10001_101010_11100;
end_screen[9][91] = 16'b10001_101010_11100;
end_screen[9][92] = 16'b10001_101010_11100;
end_screen[9][93] = 16'b10001_101010_11100;
end_screen[9][94] = 16'b10001_101010_11100;
end_screen[9][95] = 16'b10001_101010_11100;
end_screen[10][0] = 16'b10001_101010_11100;
end_screen[10][1] = 16'b10001_101010_11100;
end_screen[10][2] = 16'b10001_101010_11100;
end_screen[10][3] = 16'b10001_101010_11100;
end_screen[10][4] = 16'b10001_101010_11100;
end_screen[10][5] = 16'b10001_101010_11100;
end_screen[10][6] = 16'b10001_101010_11100;
end_screen[10][7] = 16'b10001_101010_11100;
end_screen[10][8] = 16'b10001_101010_11100;
end_screen[10][9] = 16'b10001_101010_11100;
end_screen[10][10] = 16'b10001_101010_11100;
end_screen[10][11] = 16'b10001_101010_11100;
end_screen[10][12] = 16'b10001_101010_11100;
end_screen[10][13] = 16'b10001_101010_11100;
end_screen[10][14] = 16'b10001_101010_11100;
end_screen[10][15] = 16'b10001_101010_11100;
end_screen[10][16] = 16'b10001_101010_11100;
end_screen[10][17] = 16'b10001_101010_11100;
end_screen[10][18] = 16'b01000_010100_01101;
end_screen[10][19] = 16'b00100_001000_00100;
end_screen[10][20] = 16'b00100_001000_00100;
end_screen[10][21] = 16'b00100_001000_00100;
end_screen[10][22] = 16'b00100_001000_00100;
end_screen[10][23] = 16'b00100_001000_00100;
end_screen[10][24] = 16'b00100_001000_00100;
end_screen[10][25] = 16'b00100_001000_00100;
end_screen[10][26] = 16'b01100_011101_10011;
end_screen[10][27] = 16'b10001_101010_11100;
end_screen[10][28] = 16'b10001_101010_11100;
end_screen[10][29] = 16'b01010_011001_10000;
end_screen[10][30] = 16'b00100_001000_00100;
end_screen[10][31] = 16'b00100_001000_00100;
end_screen[10][32] = 16'b00100_001000_00100;
end_screen[10][33] = 16'b01010_011001_10000;
end_screen[10][34] = 16'b10001_101010_11100;
end_screen[10][35] = 16'b10001_101010_11100;
end_screen[10][36] = 16'b00101_001011_00111;
end_screen[10][37] = 16'b00100_001000_00100;
end_screen[10][38] = 16'b00100_001000_00100;
end_screen[10][39] = 16'b00100_001000_00100;
end_screen[10][40] = 16'b00100_001000_00100;
end_screen[10][41] = 16'b00100_001000_00100;
end_screen[10][42] = 16'b00100_001000_00100;
end_screen[10][43] = 16'b00100_001000_00100;
end_screen[10][44] = 16'b00100_001000_00100;
end_screen[10][45] = 16'b00110_001111_01001;
end_screen[10][46] = 16'b10000_101000_11011;
end_screen[10][47] = 16'b10001_101010_11100;
end_screen[10][48] = 16'b10001_101010_11100;
end_screen[10][49] = 16'b00110_001111_01001;
end_screen[10][50] = 16'b00100_001000_00100;
end_screen[10][51] = 16'b00100_001000_00100;
end_screen[10][52] = 16'b00100_001000_00100;
end_screen[10][53] = 16'b01101_011111_10101;
end_screen[10][54] = 16'b10001_101010_11100;
end_screen[10][55] = 16'b10001_101010_11100;
end_screen[10][56] = 16'b01010_011001_10000;
end_screen[10][57] = 16'b00100_001000_00100;
end_screen[10][58] = 16'b00100_001000_00100;
end_screen[10][59] = 16'b00100_001000_00100;
end_screen[10][60] = 16'b00100_001000_00100;
end_screen[10][61] = 16'b00100_001000_00100;
end_screen[10][62] = 16'b00100_001000_00100;
end_screen[10][63] = 16'b00100_001000_00100;
end_screen[10][64] = 16'b01010_011001_10000;
end_screen[10][65] = 16'b10001_101010_11100;
end_screen[10][66] = 16'b10001_101010_11100;
end_screen[10][67] = 16'b00100_001000_00100;
end_screen[10][68] = 16'b00100_001000_00100;
end_screen[10][69] = 16'b00100_001000_00100;
end_screen[10][70] = 16'b00100_001000_00100;
end_screen[10][71] = 16'b00100_001000_00100;
end_screen[10][72] = 16'b00100_001000_00100;
end_screen[10][73] = 16'b00100_001000_00100;
end_screen[10][74] = 16'b00100_001000_00100;
end_screen[10][75] = 16'b00100_001000_00100;
end_screen[10][76] = 16'b00100_001000_00100;
end_screen[10][77] = 16'b01101_100001_10110;
end_screen[10][78] = 16'b10001_101010_11100;
end_screen[10][79] = 16'b10001_101010_11100;
end_screen[10][80] = 16'b10001_101010_11100;
end_screen[10][81] = 16'b10001_101010_11100;
end_screen[10][82] = 16'b10001_101010_11100;
end_screen[10][83] = 16'b10001_101010_11100;
end_screen[10][84] = 16'b10001_101010_11100;
end_screen[10][85] = 16'b10001_101010_11100;
end_screen[10][86] = 16'b10001_101010_11100;
end_screen[10][87] = 16'b10001_101010_11100;
end_screen[10][88] = 16'b10001_101010_11100;
end_screen[10][89] = 16'b10001_101010_11100;
end_screen[10][90] = 16'b10001_101010_11100;
end_screen[10][91] = 16'b10001_101010_11100;
end_screen[10][92] = 16'b10001_101010_11100;
end_screen[10][93] = 16'b10001_101010_11100;
end_screen[10][94] = 16'b10001_101010_11100;
end_screen[10][95] = 16'b10001_101010_11100;
end_screen[11][0] = 16'b10001_101010_11100;
end_screen[11][1] = 16'b10001_101010_11100;
end_screen[11][2] = 16'b10001_101010_11100;
end_screen[11][3] = 16'b10001_101010_11100;
end_screen[11][4] = 16'b10001_101010_11100;
end_screen[11][5] = 16'b10001_101010_11100;
end_screen[11][6] = 16'b10001_101010_11100;
end_screen[11][7] = 16'b10001_101010_11100;
end_screen[11][8] = 16'b10001_101010_11100;
end_screen[11][9] = 16'b10001_101010_11100;
end_screen[11][10] = 16'b10001_101010_11100;
end_screen[11][11] = 16'b10001_101010_11100;
end_screen[11][12] = 16'b10001_101010_11100;
end_screen[11][13] = 16'b10001_101010_11100;
end_screen[11][14] = 16'b10001_101010_11100;
end_screen[11][15] = 16'b10001_101010_11100;
end_screen[11][16] = 16'b10001_101010_11100;
end_screen[11][17] = 16'b10001_101010_11100;
end_screen[11][18] = 16'b01000_010100_01101;
end_screen[11][19] = 16'b00100_001000_00100;
end_screen[11][20] = 16'b00100_001000_00100;
end_screen[11][21] = 16'b00100_001000_00100;
end_screen[11][22] = 16'b00100_001000_00100;
end_screen[11][23] = 16'b00100_001000_00100;
end_screen[11][24] = 16'b00100_001000_00100;
end_screen[11][25] = 16'b00100_001000_00100;
end_screen[11][26] = 16'b00100_001000_00100;
end_screen[11][27] = 16'b10000_101000_11011;
end_screen[11][28] = 16'b10001_101010_11100;
end_screen[11][29] = 16'b01010_011001_10000;
end_screen[11][30] = 16'b00100_001000_00100;
end_screen[11][31] = 16'b00100_001000_00100;
end_screen[11][32] = 16'b00100_001000_00100;
end_screen[11][33] = 16'b01010_011001_10000;
end_screen[11][34] = 16'b10001_101010_11100;
end_screen[11][35] = 16'b10001_101010_11100;
end_screen[11][36] = 16'b00100_001000_00100;
end_screen[11][37] = 16'b00100_001000_00100;
end_screen[11][38] = 16'b00100_001000_00100;
end_screen[11][39] = 16'b00100_001000_00100;
end_screen[11][40] = 16'b00100_001000_00100;
end_screen[11][41] = 16'b00100_001000_00100;
end_screen[11][42] = 16'b00100_001000_00100;
end_screen[11][43] = 16'b00100_001000_00100;
end_screen[11][44] = 16'b00100_001000_00100;
end_screen[11][45] = 16'b00100_001000_00100;
end_screen[11][46] = 16'b01100_011101_10011;
end_screen[11][47] = 16'b10001_101010_11100;
end_screen[11][48] = 16'b10001_101010_11100;
end_screen[11][49] = 16'b00110_001111_01001;
end_screen[11][50] = 16'b00100_001000_00100;
end_screen[11][51] = 16'b00100_001000_00100;
end_screen[11][52] = 16'b00100_001000_00100;
end_screen[11][53] = 16'b01101_011111_10101;
end_screen[11][54] = 16'b10001_101010_11100;
end_screen[11][55] = 16'b10001_101010_11100;
end_screen[11][56] = 16'b00100_001000_00100;
end_screen[11][57] = 16'b00100_001000_00100;
end_screen[11][58] = 16'b00100_001000_00100;
end_screen[11][59] = 16'b00100_001000_00100;
end_screen[11][60] = 16'b01011_011011_10010;
end_screen[11][61] = 16'b01100_011101_10011;
end_screen[11][62] = 16'b01011_011011_10010;
end_screen[11][63] = 16'b01001_010111_01111;
end_screen[11][64] = 16'b01111_100101_11001;
end_screen[11][65] = 16'b10001_101010_11100;
end_screen[11][66] = 16'b10001_101010_11100;
end_screen[11][67] = 16'b00100_001000_00100;
end_screen[11][68] = 16'b00100_001000_00100;
end_screen[11][69] = 16'b00100_001000_00100;
end_screen[11][70] = 16'b00100_001000_00100;
end_screen[11][71] = 16'b00100_001000_00100;
end_screen[11][72] = 16'b00100_001000_00100;
end_screen[11][73] = 16'b00100_001000_00100;
end_screen[11][74] = 16'b00100_001000_00100;
end_screen[11][75] = 16'b00100_001000_00100;
end_screen[11][76] = 16'b00100_001000_00100;
end_screen[11][77] = 16'b01010_011001_10000;
end_screen[11][78] = 16'b10001_101010_11100;
end_screen[11][79] = 16'b10001_101010_11100;
end_screen[11][80] = 16'b10001_101010_11100;
end_screen[11][81] = 16'b10001_101010_11100;
end_screen[11][82] = 16'b10001_101010_11100;
end_screen[11][83] = 16'b10001_101010_11100;
end_screen[11][84] = 16'b10001_101010_11100;
end_screen[11][85] = 16'b10001_101010_11100;
end_screen[11][86] = 16'b10001_101010_11100;
end_screen[11][87] = 16'b10001_101010_11100;
end_screen[11][88] = 16'b10001_101010_11100;
end_screen[11][89] = 16'b10001_101010_11100;
end_screen[11][90] = 16'b10001_101010_11100;
end_screen[11][91] = 16'b10001_101010_11100;
end_screen[11][92] = 16'b10001_101010_11100;
end_screen[11][93] = 16'b10001_101010_11100;
end_screen[11][94] = 16'b10001_101010_11100;
end_screen[11][95] = 16'b10001_101010_11100;
end_screen[12][0] = 16'b10001_101010_11100;
end_screen[12][1] = 16'b10001_101010_11100;
end_screen[12][2] = 16'b10001_101010_11100;
end_screen[12][3] = 16'b10001_101010_11100;
end_screen[12][4] = 16'b10001_101010_11100;
end_screen[12][5] = 16'b10001_101010_11100;
end_screen[12][6] = 16'b10001_101010_11100;
end_screen[12][7] = 16'b10001_101010_11100;
end_screen[12][8] = 16'b10001_101010_11100;
end_screen[12][9] = 16'b10001_101010_11100;
end_screen[12][10] = 16'b10001_101010_11100;
end_screen[12][11] = 16'b10001_101010_11100;
end_screen[12][12] = 16'b10001_101010_11100;
end_screen[12][13] = 16'b10001_101010_11100;
end_screen[12][14] = 16'b10001_101010_11100;
end_screen[12][15] = 16'b10001_101010_11100;
end_screen[12][16] = 16'b10001_101010_11100;
end_screen[12][17] = 16'b10001_101010_11100;
end_screen[12][18] = 16'b01000_010100_01101;
end_screen[12][19] = 16'b00100_001000_00100;
end_screen[12][20] = 16'b00100_001000_00100;
end_screen[12][21] = 16'b00100_001000_00100;
end_screen[12][22] = 16'b00100_001000_00100;
end_screen[12][23] = 16'b00100_001000_00100;
end_screen[12][24] = 16'b00100_001000_00100;
end_screen[12][25] = 16'b00100_001000_00100;
end_screen[12][26] = 16'b00100_001000_00100;
end_screen[12][27] = 16'b10000_101000_11011;
end_screen[12][28] = 16'b10001_101010_11100;
end_screen[12][29] = 16'b01010_011001_10000;
end_screen[12][30] = 16'b00100_001000_00100;
end_screen[12][31] = 16'b00100_001000_00100;
end_screen[12][32] = 16'b00100_001000_00100;
end_screen[12][33] = 16'b01010_011001_10000;
end_screen[12][34] = 16'b10001_101010_11100;
end_screen[12][35] = 16'b10001_101010_11100;
end_screen[12][36] = 16'b00100_001000_00100;
end_screen[12][37] = 16'b00100_001000_00100;
end_screen[12][38] = 16'b00100_001000_00100;
end_screen[12][39] = 16'b00100_001000_00100;
end_screen[12][40] = 16'b01100_011101_10011;
end_screen[12][41] = 16'b10001_101010_11100;
end_screen[12][42] = 16'b00111_010001_01011;
end_screen[12][43] = 16'b00100_001000_00100;
end_screen[12][44] = 16'b00100_001000_00100;
end_screen[12][45] = 16'b00100_001000_00100;
end_screen[12][46] = 16'b01010_011001_10000;
end_screen[12][47] = 16'b10001_101010_11100;
end_screen[12][48] = 16'b10001_101010_11100;
end_screen[12][49] = 16'b00110_001111_01001;
end_screen[12][50] = 16'b00100_001000_00100;
end_screen[12][51] = 16'b00100_001000_00100;
end_screen[12][52] = 16'b00100_001000_00100;
end_screen[12][53] = 16'b01101_011111_10101;
end_screen[12][54] = 16'b10001_101010_11100;
end_screen[12][55] = 16'b10001_101010_11100;
end_screen[12][56] = 16'b00111_010001_01011;
end_screen[12][57] = 16'b00100_001000_00100;
end_screen[12][58] = 16'b00100_001000_00100;
end_screen[12][59] = 16'b00100_001000_00100;
end_screen[12][60] = 16'b00100_001000_00100;
end_screen[12][61] = 16'b01001_010111_01111;
end_screen[12][62] = 16'b01100_011101_10011;
end_screen[12][63] = 16'b10001_101010_11100;
end_screen[12][64] = 16'b10001_101010_11100;
end_screen[12][65] = 16'b10001_101010_11100;
end_screen[12][66] = 16'b10001_101010_11100;
end_screen[12][67] = 16'b00100_001000_00100;
end_screen[12][68] = 16'b00100_001000_00100;
end_screen[12][69] = 16'b00100_001000_00100;
end_screen[12][70] = 16'b00100_001000_00100;
end_screen[12][71] = 16'b01101_011111_10101;
end_screen[12][72] = 16'b10001_101010_11100;
end_screen[12][73] = 16'b01000_010100_01101;
end_screen[12][74] = 16'b00100_001000_00100;
end_screen[12][75] = 16'b00100_001000_00100;
end_screen[12][76] = 16'b00100_001000_00100;
end_screen[12][77] = 16'b01010_011001_10000;
end_screen[12][78] = 16'b10001_101010_11100;
end_screen[12][79] = 16'b10001_101010_11100;
end_screen[12][80] = 16'b10001_101010_11100;
end_screen[12][81] = 16'b10001_101010_11100;
end_screen[12][82] = 16'b10001_101010_11100;
end_screen[12][83] = 16'b10001_101010_11100;
end_screen[12][84] = 16'b10001_101010_11100;
end_screen[12][85] = 16'b10001_101010_11100;
end_screen[12][86] = 16'b10001_101010_11100;
end_screen[12][87] = 16'b10001_101010_11100;
end_screen[12][88] = 16'b10001_101010_11100;
end_screen[12][89] = 16'b10001_101010_11100;
end_screen[12][90] = 16'b10001_101010_11100;
end_screen[12][91] = 16'b10001_101010_11100;
end_screen[12][92] = 16'b10001_101010_11100;
end_screen[12][93] = 16'b10001_101010_11100;
end_screen[12][94] = 16'b10001_101010_11100;
end_screen[12][95] = 16'b10001_101010_11100;
end_screen[13][0] = 16'b10001_101010_11100;
end_screen[13][1] = 16'b10001_101010_11100;
end_screen[13][2] = 16'b10001_101010_11100;
end_screen[13][3] = 16'b10001_101010_11100;
end_screen[13][4] = 16'b10001_101010_11100;
end_screen[13][5] = 16'b10001_101010_11100;
end_screen[13][6] = 16'b10001_101010_11100;
end_screen[13][7] = 16'b10001_101010_11100;
end_screen[13][8] = 16'b10001_101010_11100;
end_screen[13][9] = 16'b10001_101010_11100;
end_screen[13][10] = 16'b10001_101010_11100;
end_screen[13][11] = 16'b10001_101010_11100;
end_screen[13][12] = 16'b10001_101010_11100;
end_screen[13][13] = 16'b10001_101010_11100;
end_screen[13][14] = 16'b10001_101010_11100;
end_screen[13][15] = 16'b10001_101010_11100;
end_screen[13][16] = 16'b10001_101010_11100;
end_screen[13][17] = 16'b10001_101010_11100;
end_screen[13][18] = 16'b01000_010100_01101;
end_screen[13][19] = 16'b00100_001000_00100;
end_screen[13][20] = 16'b00100_001000_00100;
end_screen[13][21] = 16'b00100_001000_00100;
end_screen[13][22] = 16'b00100_001000_00100;
end_screen[13][23] = 16'b00100_001000_00100;
end_screen[13][24] = 16'b00100_001000_00100;
end_screen[13][25] = 16'b00100_001000_00100;
end_screen[13][26] = 16'b01101_011111_10101;
end_screen[13][27] = 16'b10001_101010_11100;
end_screen[13][28] = 16'b10001_101010_11100;
end_screen[13][29] = 16'b01010_011001_10000;
end_screen[13][30] = 16'b00100_001000_00100;
end_screen[13][31] = 16'b00100_001000_00100;
end_screen[13][32] = 16'b00100_001000_00100;
end_screen[13][33] = 16'b01010_011001_10000;
end_screen[13][34] = 16'b10001_101010_11100;
end_screen[13][35] = 16'b10001_101010_11100;
end_screen[13][36] = 16'b00100_001000_00100;
end_screen[13][37] = 16'b00100_001000_00100;
end_screen[13][38] = 16'b00100_001000_00100;
end_screen[13][39] = 16'b00100_001000_00100;
end_screen[13][40] = 16'b01110_100011_10111;
end_screen[13][41] = 16'b10001_101010_11100;
end_screen[13][42] = 16'b01010_011001_10000;
end_screen[13][43] = 16'b00100_001000_00100;
end_screen[13][44] = 16'b00100_001000_00100;
end_screen[13][45] = 16'b00100_001000_00100;
end_screen[13][46] = 16'b01010_011001_10000;
end_screen[13][47] = 16'b10001_101010_11100;
end_screen[13][48] = 16'b10001_101010_11100;
end_screen[13][49] = 16'b00110_001111_01001;
end_screen[13][50] = 16'b00100_001000_00100;
end_screen[13][51] = 16'b00100_001000_00100;
end_screen[13][52] = 16'b00100_001000_00100;
end_screen[13][53] = 16'b01101_011111_10101;
end_screen[13][54] = 16'b10001_101010_11100;
end_screen[13][55] = 16'b10001_101010_11100;
end_screen[13][56] = 16'b01101_100001_10110;
end_screen[13][57] = 16'b00100_001000_00100;
end_screen[13][58] = 16'b00100_001000_00100;
end_screen[13][59] = 16'b00100_001000_00100;
end_screen[13][60] = 16'b00100_001000_00100;
end_screen[13][61] = 16'b00100_001000_00100;
end_screen[13][62] = 16'b00100_001000_00100;
end_screen[13][63] = 16'b00110_001111_01001;
end_screen[13][64] = 16'b10000_100111_11010;
end_screen[13][65] = 16'b10001_101010_11100;
end_screen[13][66] = 16'b10001_101010_11100;
end_screen[13][67] = 16'b00100_001000_00100;
end_screen[13][68] = 16'b00100_001000_00100;
end_screen[13][69] = 16'b00100_001000_00100;
end_screen[13][70] = 16'b00100_001000_00100;
end_screen[13][71] = 16'b01110_100011_10111;
end_screen[13][72] = 16'b10001_101010_11100;
end_screen[13][73] = 16'b01010_011001_10000;
end_screen[13][74] = 16'b00100_001000_00100;
end_screen[13][75] = 16'b00100_001000_00100;
end_screen[13][76] = 16'b00100_001000_00100;
end_screen[13][77] = 16'b01010_011001_10000;
end_screen[13][78] = 16'b10001_101010_11100;
end_screen[13][79] = 16'b10001_101010_11100;
end_screen[13][80] = 16'b10001_101010_11100;
end_screen[13][81] = 16'b10001_101010_11100;
end_screen[13][82] = 16'b10001_101010_11100;
end_screen[13][83] = 16'b10001_101010_11100;
end_screen[13][84] = 16'b10001_101010_11100;
end_screen[13][85] = 16'b10001_101010_11100;
end_screen[13][86] = 16'b10001_101010_11100;
end_screen[13][87] = 16'b10001_101010_11100;
end_screen[13][88] = 16'b10001_101010_11100;
end_screen[13][89] = 16'b10001_101010_11100;
end_screen[13][90] = 16'b10001_101010_11100;
end_screen[13][91] = 16'b10001_101010_11100;
end_screen[13][92] = 16'b10001_101010_11100;
end_screen[13][93] = 16'b10001_101010_11100;
end_screen[13][94] = 16'b10001_101010_11100;
end_screen[13][95] = 16'b10001_101010_11100;
end_screen[14][0] = 16'b10001_101010_11100;
end_screen[14][1] = 16'b10001_101010_11100;
end_screen[14][2] = 16'b10001_101010_11100;
end_screen[14][3] = 16'b10001_101010_11100;
end_screen[14][4] = 16'b10001_101010_11100;
end_screen[14][5] = 16'b10001_101010_11100;
end_screen[14][6] = 16'b10001_101010_11100;
end_screen[14][7] = 16'b10001_101010_11100;
end_screen[14][8] = 16'b10001_101010_11100;
end_screen[14][9] = 16'b10001_101010_11100;
end_screen[14][10] = 16'b10001_101010_11100;
end_screen[14][11] = 16'b10001_101010_11100;
end_screen[14][12] = 16'b10001_101010_11100;
end_screen[14][13] = 16'b10001_101010_11100;
end_screen[14][14] = 16'b10001_101010_11100;
end_screen[14][15] = 16'b10001_101010_11100;
end_screen[14][16] = 16'b10001_101010_11100;
end_screen[14][17] = 16'b10001_101010_11100;
end_screen[14][18] = 16'b01000_010100_01101;
end_screen[14][19] = 16'b00100_001000_00100;
end_screen[14][20] = 16'b00100_001000_00100;
end_screen[14][21] = 16'b00100_001000_00100;
end_screen[14][22] = 16'b01000_010100_01101;
end_screen[14][23] = 16'b10001_101010_11100;
end_screen[14][24] = 16'b10001_101010_11100;
end_screen[14][25] = 16'b10001_101010_11100;
end_screen[14][26] = 16'b10001_101010_11100;
end_screen[14][27] = 16'b10001_101010_11100;
end_screen[14][28] = 16'b10001_101010_11100;
end_screen[14][29] = 16'b01010_011001_10000;
end_screen[14][30] = 16'b00100_001000_00100;
end_screen[14][31] = 16'b00100_001000_00100;
end_screen[14][32] = 16'b00100_001000_00100;
end_screen[14][33] = 16'b01010_011001_10000;
end_screen[14][34] = 16'b10001_101010_11100;
end_screen[14][35] = 16'b10001_101010_11100;
end_screen[14][36] = 16'b00100_001000_00100;
end_screen[14][37] = 16'b00100_001000_00100;
end_screen[14][38] = 16'b00100_001000_00100;
end_screen[14][39] = 16'b00100_001000_00100;
end_screen[14][40] = 16'b01110_100011_10111;
end_screen[14][41] = 16'b10001_101010_11100;
end_screen[14][42] = 16'b01010_011001_10000;
end_screen[14][43] = 16'b00100_001000_00100;
end_screen[14][44] = 16'b00100_001000_00100;
end_screen[14][45] = 16'b00100_001000_00100;
end_screen[14][46] = 16'b01010_011001_10000;
end_screen[14][47] = 16'b10001_101010_11100;
end_screen[14][48] = 16'b10001_101010_11100;
end_screen[14][49] = 16'b00110_001111_01001;
end_screen[14][50] = 16'b00100_001000_00100;
end_screen[14][51] = 16'b00100_001000_00100;
end_screen[14][52] = 16'b00100_001000_00100;
end_screen[14][53] = 16'b01101_011111_10101;
end_screen[14][54] = 16'b10001_101010_11100;
end_screen[14][55] = 16'b10001_101010_11100;
end_screen[14][56] = 16'b10001_101010_11100;
end_screen[14][57] = 16'b01111_100101_11001;
end_screen[14][58] = 16'b01100_011101_10011;
end_screen[14][59] = 16'b00101_001011_00111;
end_screen[14][60] = 16'b00100_001000_00100;
end_screen[14][61] = 16'b00100_001000_00100;
end_screen[14][62] = 16'b00100_001000_00100;
end_screen[14][63] = 16'b00100_001000_00100;
end_screen[14][64] = 16'b01001_010111_01111;
end_screen[14][65] = 16'b10001_101010_11100;
end_screen[14][66] = 16'b10001_101010_11100;
end_screen[14][67] = 16'b00100_001000_00100;
end_screen[14][68] = 16'b00100_001000_00100;
end_screen[14][69] = 16'b00100_001000_00100;
end_screen[14][70] = 16'b00100_001000_00100;
end_screen[14][71] = 16'b01110_100011_10111;
end_screen[14][72] = 16'b10001_101010_11100;
end_screen[14][73] = 16'b01010_011001_10000;
end_screen[14][74] = 16'b00100_001000_00100;
end_screen[14][75] = 16'b00100_001000_00100;
end_screen[14][76] = 16'b00100_001000_00100;
end_screen[14][77] = 16'b01010_011001_10000;
end_screen[14][78] = 16'b10001_101010_11100;
end_screen[14][79] = 16'b10001_101010_11100;
end_screen[14][80] = 16'b10001_101010_11100;
end_screen[14][81] = 16'b10001_101010_11100;
end_screen[14][82] = 16'b10001_101010_11100;
end_screen[14][83] = 16'b10001_101010_11100;
end_screen[14][84] = 16'b10001_101010_11100;
end_screen[14][85] = 16'b10001_101010_11100;
end_screen[14][86] = 16'b10001_101010_11100;
end_screen[14][87] = 16'b10001_101010_11100;
end_screen[14][88] = 16'b10001_101010_11100;
end_screen[14][89] = 16'b10001_101010_11100;
end_screen[14][90] = 16'b10001_101010_11100;
end_screen[14][91] = 16'b10001_101010_11100;
end_screen[14][92] = 16'b10001_101010_11100;
end_screen[14][93] = 16'b10001_101010_11100;
end_screen[14][94] = 16'b10001_101010_11100;
end_screen[14][95] = 16'b10001_101010_11100;
end_screen[15][0] = 16'b10001_101010_11100;
end_screen[15][1] = 16'b10001_101010_11100;
end_screen[15][2] = 16'b10001_101010_11100;
end_screen[15][3] = 16'b10001_101010_11100;
end_screen[15][4] = 16'b10001_101010_11100;
end_screen[15][5] = 16'b10001_101010_11100;
end_screen[15][6] = 16'b10001_101010_11100;
end_screen[15][7] = 16'b10001_101010_11100;
end_screen[15][8] = 16'b10001_101010_11100;
end_screen[15][9] = 16'b10001_101010_11100;
end_screen[15][10] = 16'b10001_101010_11100;
end_screen[15][11] = 16'b10001_101010_11100;
end_screen[15][12] = 16'b10001_101010_11100;
end_screen[15][13] = 16'b10001_101010_11100;
end_screen[15][14] = 16'b10001_101010_11100;
end_screen[15][15] = 16'b10001_101010_11100;
end_screen[15][16] = 16'b10001_101010_11100;
end_screen[15][17] = 16'b10001_101010_11100;
end_screen[15][18] = 16'b01000_010100_01101;
end_screen[15][19] = 16'b00100_001000_00100;
end_screen[15][20] = 16'b00100_001000_00100;
end_screen[15][21] = 16'b00100_001000_00100;
end_screen[15][22] = 16'b01000_010100_01101;
end_screen[15][23] = 16'b10001_101010_11100;
end_screen[15][24] = 16'b10001_101010_11100;
end_screen[15][25] = 16'b10001_101010_11100;
end_screen[15][26] = 16'b10001_101010_11100;
end_screen[15][27] = 16'b10001_101010_11100;
end_screen[15][28] = 16'b10001_101010_11100;
end_screen[15][29] = 16'b01010_011001_10000;
end_screen[15][30] = 16'b00100_001000_00100;
end_screen[15][31] = 16'b00100_001000_00100;
end_screen[15][32] = 16'b00100_001000_00100;
end_screen[15][33] = 16'b01010_011001_10000;
end_screen[15][34] = 16'b10001_101010_11100;
end_screen[15][35] = 16'b10001_101010_11100;
end_screen[15][36] = 16'b00100_001000_00100;
end_screen[15][37] = 16'b00100_001000_00100;
end_screen[15][38] = 16'b00100_001000_00100;
end_screen[15][39] = 16'b00100_001000_00100;
end_screen[15][40] = 16'b01110_100011_10111;
end_screen[15][41] = 16'b10001_101010_11100;
end_screen[15][42] = 16'b01010_011001_10000;
end_screen[15][43] = 16'b00100_001000_00100;
end_screen[15][44] = 16'b00100_001000_00100;
end_screen[15][45] = 16'b00100_001000_00100;
end_screen[15][46] = 16'b01010_011001_10000;
end_screen[15][47] = 16'b10001_101010_11100;
end_screen[15][48] = 16'b10001_101010_11100;
end_screen[15][49] = 16'b00110_001111_01001;
end_screen[15][50] = 16'b00100_001000_00100;
end_screen[15][51] = 16'b00100_001000_00100;
end_screen[15][52] = 16'b00100_001000_00100;
end_screen[15][53] = 16'b01101_011111_10101;
end_screen[15][54] = 16'b10001_101010_11100;
end_screen[15][55] = 16'b10001_101010_11100;
end_screen[15][56] = 16'b01001_010111_01111;
end_screen[15][57] = 16'b00100_001000_00100;
end_screen[15][58] = 16'b01010_011001_10000;
end_screen[15][59] = 16'b01100_011101_10011;
end_screen[15][60] = 16'b01101_011111_10101;
end_screen[15][61] = 16'b00100_001000_00100;
end_screen[15][62] = 16'b00100_001000_00100;
end_screen[15][63] = 16'b00100_001000_00100;
end_screen[15][64] = 16'b00110_001111_01001;
end_screen[15][65] = 16'b10001_101010_11100;
end_screen[15][66] = 16'b10001_101010_11100;
end_screen[15][67] = 16'b00100_001000_00100;
end_screen[15][68] = 16'b00100_001000_00100;
end_screen[15][69] = 16'b00100_001000_00100;
end_screen[15][70] = 16'b00100_001000_00100;
end_screen[15][71] = 16'b01110_100011_10111;
end_screen[15][72] = 16'b10001_101010_11100;
end_screen[15][73] = 16'b01010_011001_10000;
end_screen[15][74] = 16'b00100_001000_00100;
end_screen[15][75] = 16'b00100_001000_00100;
end_screen[15][76] = 16'b00100_001000_00100;
end_screen[15][77] = 16'b01010_011001_10000;
end_screen[15][78] = 16'b10001_101010_11100;
end_screen[15][79] = 16'b10001_101010_11100;
end_screen[15][80] = 16'b10001_101010_11100;
end_screen[15][81] = 16'b10001_101010_11100;
end_screen[15][82] = 16'b10001_101010_11100;
end_screen[15][83] = 16'b10001_101010_11100;
end_screen[15][84] = 16'b10001_101010_11100;
end_screen[15][85] = 16'b10001_101010_11100;
end_screen[15][86] = 16'b10001_101010_11100;
end_screen[15][87] = 16'b10001_101010_11100;
end_screen[15][88] = 16'b10001_101010_11100;
end_screen[15][89] = 16'b10001_101010_11100;
end_screen[15][90] = 16'b10001_101010_11100;
end_screen[15][91] = 16'b10001_101010_11100;
end_screen[15][92] = 16'b10001_101010_11100;
end_screen[15][93] = 16'b10001_101010_11100;
end_screen[15][94] = 16'b10001_101010_11100;
end_screen[15][95] = 16'b10001_101010_11100;
end_screen[16][0] = 16'b10001_101010_11100;
end_screen[16][1] = 16'b10001_101010_11100;
end_screen[16][2] = 16'b10001_101010_11100;
end_screen[16][3] = 16'b10001_101010_11100;
end_screen[16][4] = 16'b10001_101010_11100;
end_screen[16][5] = 16'b10001_101010_11100;
end_screen[16][6] = 16'b10001_101010_11100;
end_screen[16][7] = 16'b10001_101010_11100;
end_screen[16][8] = 16'b10001_101010_11100;
end_screen[16][9] = 16'b10001_101010_11100;
end_screen[16][10] = 16'b10001_101010_11100;
end_screen[16][11] = 16'b10001_101010_11100;
end_screen[16][12] = 16'b10001_101010_11100;
end_screen[16][13] = 16'b10001_101010_11100;
end_screen[16][14] = 16'b10001_101010_11100;
end_screen[16][15] = 16'b10001_101010_11100;
end_screen[16][16] = 16'b10001_101010_11100;
end_screen[16][17] = 16'b10001_101010_11100;
end_screen[16][18] = 16'b01000_010100_01101;
end_screen[16][19] = 16'b00100_001000_00100;
end_screen[16][20] = 16'b00100_001000_00100;
end_screen[16][21] = 16'b00100_001000_00100;
end_screen[16][22] = 16'b01000_010100_01101;
end_screen[16][23] = 16'b10001_101010_11100;
end_screen[16][24] = 16'b10001_101010_11100;
end_screen[16][25] = 16'b10001_101010_11100;
end_screen[16][26] = 16'b10001_101010_11100;
end_screen[16][27] = 16'b10001_101010_11100;
end_screen[16][28] = 16'b10001_101010_11100;
end_screen[16][29] = 16'b01010_011001_10000;
end_screen[16][30] = 16'b00100_001000_00100;
end_screen[16][31] = 16'b00100_001000_00100;
end_screen[16][32] = 16'b00100_001000_00100;
end_screen[16][33] = 16'b01010_011001_10000;
end_screen[16][34] = 16'b10001_101010_11100;
end_screen[16][35] = 16'b10001_101010_11100;
end_screen[16][36] = 16'b00100_001000_00100;
end_screen[16][37] = 16'b00100_001000_00100;
end_screen[16][38] = 16'b00100_001000_00100;
end_screen[16][39] = 16'b00100_001000_00100;
end_screen[16][40] = 16'b01110_100011_10111;
end_screen[16][41] = 16'b10001_101010_11100;
end_screen[16][42] = 16'b01010_011001_10000;
end_screen[16][43] = 16'b00100_001000_00100;
end_screen[16][44] = 16'b00100_001000_00100;
end_screen[16][45] = 16'b00100_001000_00100;
end_screen[16][46] = 16'b01010_011001_10000;
end_screen[16][47] = 16'b10001_101010_11100;
end_screen[16][48] = 16'b10001_101010_11100;
end_screen[16][49] = 16'b00110_001111_01001;
end_screen[16][50] = 16'b00100_001000_00100;
end_screen[16][51] = 16'b00100_001000_00100;
end_screen[16][52] = 16'b00100_001000_00100;
end_screen[16][53] = 16'b01101_011111_10101;
end_screen[16][54] = 16'b10001_101010_11100;
end_screen[16][55] = 16'b01101_100001_10110;
end_screen[16][56] = 16'b00100_001000_00100;
end_screen[16][57] = 16'b00100_001000_00100;
end_screen[16][58] = 16'b00100_001000_00100;
end_screen[16][59] = 16'b00100_001000_00100;
end_screen[16][60] = 16'b00100_001000_00100;
end_screen[16][61] = 16'b00100_001000_00100;
end_screen[16][62] = 16'b00100_001000_00100;
end_screen[16][63] = 16'b00100_001000_00100;
end_screen[16][64] = 16'b00111_010001_01011;
end_screen[16][65] = 16'b10001_101010_11100;
end_screen[16][66] = 16'b10001_101010_11100;
end_screen[16][67] = 16'b00100_001000_00100;
end_screen[16][68] = 16'b00100_001000_00100;
end_screen[16][69] = 16'b00100_001000_00100;
end_screen[16][70] = 16'b00100_001000_00100;
end_screen[16][71] = 16'b01110_100011_10111;
end_screen[16][72] = 16'b10001_101010_11100;
end_screen[16][73] = 16'b01010_011001_10000;
end_screen[16][74] = 16'b00100_001000_00100;
end_screen[16][75] = 16'b00100_001000_00100;
end_screen[16][76] = 16'b00100_001000_00100;
end_screen[16][77] = 16'b01010_011001_10000;
end_screen[16][78] = 16'b10001_101010_11100;
end_screen[16][79] = 16'b10001_101010_11100;
end_screen[16][80] = 16'b10001_101010_11100;
end_screen[16][81] = 16'b10001_101010_11100;
end_screen[16][82] = 16'b10001_101010_11100;
end_screen[16][83] = 16'b10001_101010_11100;
end_screen[16][84] = 16'b10001_101010_11100;
end_screen[16][85] = 16'b10001_101010_11100;
end_screen[16][86] = 16'b10001_101010_11100;
end_screen[16][87] = 16'b10001_101010_11100;
end_screen[16][88] = 16'b10001_101010_11100;
end_screen[16][89] = 16'b10001_101010_11100;
end_screen[16][90] = 16'b10001_101010_11100;
end_screen[16][91] = 16'b10001_101010_11100;
end_screen[16][92] = 16'b10001_101010_11100;
end_screen[16][93] = 16'b10001_101010_11100;
end_screen[16][94] = 16'b10001_101010_11100;
end_screen[16][95] = 16'b10001_101010_11100;
end_screen[17][0] = 16'b10001_101010_11100;
end_screen[17][1] = 16'b10001_101010_11100;
end_screen[17][2] = 16'b10001_101010_11100;
end_screen[17][3] = 16'b10001_101010_11100;
end_screen[17][4] = 16'b10001_101010_11100;
end_screen[17][5] = 16'b10001_101010_11100;
end_screen[17][6] = 16'b10001_101010_11100;
end_screen[17][7] = 16'b10001_101010_11100;
end_screen[17][8] = 16'b10001_101010_11100;
end_screen[17][9] = 16'b10001_101010_11100;
end_screen[17][10] = 16'b10001_101010_11100;
end_screen[17][11] = 16'b10001_101010_11100;
end_screen[17][12] = 16'b10001_101010_11100;
end_screen[17][13] = 16'b10001_101010_11100;
end_screen[17][14] = 16'b10001_101010_11100;
end_screen[17][15] = 16'b10001_101010_11100;
end_screen[17][16] = 16'b10001_101010_11100;
end_screen[17][17] = 16'b10001_101010_11100;
end_screen[17][18] = 16'b01011_011011_10010;
end_screen[17][19] = 16'b00100_001000_00100;
end_screen[17][20] = 16'b00100_001000_00100;
end_screen[17][21] = 16'b00100_001000_00100;
end_screen[17][22] = 16'b01011_011011_10010;
end_screen[17][23] = 16'b10001_101010_11100;
end_screen[17][24] = 16'b10001_101010_11100;
end_screen[17][25] = 16'b10001_101010_11100;
end_screen[17][26] = 16'b10001_101010_11100;
end_screen[17][27] = 16'b10001_101010_11100;
end_screen[17][28] = 16'b10001_101010_11100;
end_screen[17][29] = 16'b01011_011011_10010;
end_screen[17][30] = 16'b00100_001000_00100;
end_screen[17][31] = 16'b00100_001000_00100;
end_screen[17][32] = 16'b00100_001000_00100;
end_screen[17][33] = 16'b01100_011101_10011;
end_screen[17][34] = 16'b10001_101010_11100;
end_screen[17][35] = 16'b10001_101010_11100;
end_screen[17][36] = 16'b00101_001011_00111;
end_screen[17][37] = 16'b00100_001000_00100;
end_screen[17][38] = 16'b00100_001000_00100;
end_screen[17][39] = 16'b00100_001000_00100;
end_screen[17][40] = 16'b01111_100101_11001;
end_screen[17][41] = 16'b10001_101010_11100;
end_screen[17][42] = 16'b01011_011011_10010;
end_screen[17][43] = 16'b00100_001000_00100;
end_screen[17][44] = 16'b00100_001000_00100;
end_screen[17][45] = 16'b00100_001000_00100;
end_screen[17][46] = 16'b01011_011011_10010;
end_screen[17][47] = 16'b10001_101010_11100;
end_screen[17][48] = 16'b10001_101010_11100;
end_screen[17][49] = 16'b00111_010001_01011;
end_screen[17][50] = 16'b00100_001000_00100;
end_screen[17][51] = 16'b00100_001000_00100;
end_screen[17][52] = 16'b00100_001000_00100;
end_screen[17][53] = 16'b01111_100101_11001;
end_screen[17][54] = 16'b10001_101010_11100;
end_screen[17][55] = 16'b10000_101000_11011;
end_screen[17][56] = 16'b00110_001111_01001;
end_screen[17][57] = 16'b00100_001000_00100;
end_screen[17][58] = 16'b00100_001000_00100;
end_screen[17][59] = 16'b00100_001000_00100;
end_screen[17][60] = 16'b00100_001000_00100;
end_screen[17][61] = 16'b00100_001000_00100;
end_screen[17][62] = 16'b00100_001000_00100;
end_screen[17][63] = 16'b00100_001000_00100;
end_screen[17][64] = 16'b01111_100101_11001;
end_screen[17][65] = 16'b10001_101010_11100;
end_screen[17][66] = 16'b10001_101010_11100;
end_screen[17][67] = 16'b00101_001011_00111;
end_screen[17][68] = 16'b00100_001000_00100;
end_screen[17][69] = 16'b00100_001000_00100;
end_screen[17][70] = 16'b00100_001000_00100;
end_screen[17][71] = 16'b01111_100101_11001;
end_screen[17][72] = 16'b10001_101010_11100;
end_screen[17][73] = 16'b01011_011011_10010;
end_screen[17][74] = 16'b00100_001000_00100;
end_screen[17][75] = 16'b00100_001000_00100;
end_screen[17][76] = 16'b00100_001000_00100;
end_screen[17][77] = 16'b01011_011011_10010;
end_screen[17][78] = 16'b10001_101010_11100;
end_screen[17][79] = 16'b10001_101010_11100;
end_screen[17][80] = 16'b10001_101010_11100;
end_screen[17][81] = 16'b10001_101010_11100;
end_screen[17][82] = 16'b10001_101010_11100;
end_screen[17][83] = 16'b10001_101010_11100;
end_screen[17][84] = 16'b10001_101010_11100;
end_screen[17][85] = 16'b10001_101010_11100;
end_screen[17][86] = 16'b10001_101010_11100;
end_screen[17][87] = 16'b10001_101010_11100;
end_screen[17][88] = 16'b10001_101010_11100;
end_screen[17][89] = 16'b10001_101010_11100;
end_screen[17][90] = 16'b10001_101010_11100;
end_screen[17][91] = 16'b10001_101010_11100;
end_screen[17][92] = 16'b10001_101010_11100;
end_screen[17][93] = 16'b10001_101010_11100;
end_screen[17][94] = 16'b10001_101010_11100;
end_screen[17][95] = 16'b10001_101010_11100;
end_screen[18][0] = 16'b10001_101010_11100;
end_screen[18][1] = 16'b10001_101010_11100;
end_screen[18][2] = 16'b10001_101010_11100;
end_screen[18][3] = 16'b10001_101010_11100;
end_screen[18][4] = 16'b10001_101010_11100;
end_screen[18][5] = 16'b10001_101010_11100;
end_screen[18][6] = 16'b10001_101010_11100;
end_screen[18][7] = 16'b10001_101010_11100;
end_screen[18][8] = 16'b10001_101010_11100;
end_screen[18][9] = 16'b10001_101010_11100;
end_screen[18][10] = 16'b10001_101010_11100;
end_screen[18][11] = 16'b10001_101010_11100;
end_screen[18][12] = 16'b10001_101010_11100;
end_screen[18][13] = 16'b10001_101010_11100;
end_screen[18][14] = 16'b10001_101010_11100;
end_screen[18][15] = 16'b10001_101010_11100;
end_screen[18][16] = 16'b10001_101010_11100;
end_screen[18][17] = 16'b10001_101010_11100;
end_screen[18][18] = 16'b10000_101000_11011;
end_screen[18][19] = 16'b01000_010100_01101;
end_screen[18][20] = 16'b00100_001000_00100;
end_screen[18][21] = 16'b01000_010100_01101;
end_screen[18][22] = 16'b10000_101000_11011;
end_screen[18][23] = 16'b10001_101010_11100;
end_screen[18][24] = 16'b10001_101010_11100;
end_screen[18][25] = 16'b10001_101010_11100;
end_screen[18][26] = 16'b10001_101010_11100;
end_screen[18][27] = 16'b10001_101010_11100;
end_screen[18][28] = 16'b10001_101010_11100;
end_screen[18][29] = 16'b10000_101000_11011;
end_screen[18][30] = 16'b01000_010100_01101;
end_screen[18][31] = 16'b00100_001000_00100;
end_screen[18][32] = 16'b01000_010100_01101;
end_screen[18][33] = 16'b10000_101000_11011;
end_screen[18][34] = 16'b10001_101010_11100;
end_screen[18][35] = 16'b10001_101010_11100;
end_screen[18][36] = 16'b01110_100011_10111;
end_screen[18][37] = 16'b00101_001011_00111;
end_screen[18][38] = 16'b00100_001000_00100;
end_screen[18][39] = 16'b01100_011101_10011;
end_screen[18][40] = 16'b10001_101010_11100;
end_screen[18][41] = 16'b10001_101010_11100;
end_screen[18][42] = 16'b10000_101000_11011;
end_screen[18][43] = 16'b01000_010100_01101;
end_screen[18][44] = 16'b00100_001000_00100;
end_screen[18][45] = 16'b01000_010100_01101;
end_screen[18][46] = 16'b10000_101000_11011;
end_screen[18][47] = 16'b10001_101010_11100;
end_screen[18][48] = 16'b10001_101010_11100;
end_screen[18][49] = 16'b01111_100101_11001;
end_screen[18][50] = 16'b00110_001111_01001;
end_screen[18][51] = 16'b00100_001000_00100;
end_screen[18][52] = 16'b01011_011011_10010;
end_screen[18][53] = 16'b10001_101010_11100;
end_screen[18][54] = 16'b10001_101010_11100;
end_screen[18][55] = 16'b10001_101010_11100;
end_screen[18][56] = 16'b10000_101000_11011;
end_screen[18][57] = 16'b01100_011101_10011;
end_screen[18][58] = 16'b00100_001000_00100;
end_screen[18][59] = 16'b00100_001000_00100;
end_screen[18][60] = 16'b00100_001000_00100;
end_screen[18][61] = 16'b00100_001000_00100;
end_screen[18][62] = 16'b01010_011001_10000;
end_screen[18][63] = 16'b01111_100101_11001;
end_screen[18][64] = 16'b10001_101010_11100;
end_screen[18][65] = 16'b10001_101010_11100;
end_screen[18][66] = 16'b10001_101010_11100;
end_screen[18][67] = 16'b01110_100011_10111;
end_screen[18][68] = 16'b00101_001011_00111;
end_screen[18][69] = 16'b00100_001000_00100;
end_screen[18][70] = 16'b01100_011101_10011;
end_screen[18][71] = 16'b10001_101010_11100;
end_screen[18][72] = 16'b10001_101010_11100;
end_screen[18][73] = 16'b10000_101000_11011;
end_screen[18][74] = 16'b01000_010100_01101;
end_screen[18][75] = 16'b00100_001000_00100;
end_screen[18][76] = 16'b01000_010100_01101;
end_screen[18][77] = 16'b10000_101000_11011;
end_screen[18][78] = 16'b10001_101010_11100;
end_screen[18][79] = 16'b10001_101010_11100;
end_screen[18][80] = 16'b10001_101010_11100;
end_screen[18][81] = 16'b10001_101010_11100;
end_screen[18][82] = 16'b10001_101010_11100;
end_screen[18][83] = 16'b10001_101010_11100;
end_screen[18][84] = 16'b10001_101010_11100;
end_screen[18][85] = 16'b10001_101010_11100;
end_screen[18][86] = 16'b10001_101010_11100;
end_screen[18][87] = 16'b10001_101010_11100;
end_screen[18][88] = 16'b10001_101010_11100;
end_screen[18][89] = 16'b10001_101010_11100;
end_screen[18][90] = 16'b10001_101010_11100;
end_screen[18][91] = 16'b10001_101010_11100;
end_screen[18][92] = 16'b10001_101010_11100;
end_screen[18][93] = 16'b10001_101010_11100;
end_screen[18][94] = 16'b10001_101010_11100;
end_screen[18][95] = 16'b10001_101010_11100;
end_screen[19][0] = 16'b10001_101010_11100;
end_screen[19][1] = 16'b10001_101010_11100;
end_screen[19][2] = 16'b10001_101010_11100;
end_screen[19][3] = 16'b10001_101010_11100;
end_screen[19][4] = 16'b10001_101010_11100;
end_screen[19][5] = 16'b10001_101010_11100;
end_screen[19][6] = 16'b10001_101010_11100;
end_screen[19][7] = 16'b10001_101010_11100;
end_screen[19][8] = 16'b10001_101010_11100;
end_screen[19][9] = 16'b10001_101010_11100;
end_screen[19][10] = 16'b10001_101010_11100;
end_screen[19][11] = 16'b10001_101010_11100;
end_screen[19][12] = 16'b10001_101010_11100;
end_screen[19][13] = 16'b10001_101010_11100;
end_screen[19][14] = 16'b10001_101010_11100;
end_screen[19][15] = 16'b10001_101010_11100;
end_screen[19][16] = 16'b10001_101010_11100;
end_screen[19][17] = 16'b10001_101010_11100;
end_screen[19][18] = 16'b10001_101010_11100;
end_screen[19][19] = 16'b10001_101010_11100;
end_screen[19][20] = 16'b10001_101010_11100;
end_screen[19][21] = 16'b10001_101010_11100;
end_screen[19][22] = 16'b10001_101010_11100;
end_screen[19][23] = 16'b10001_101010_11100;
end_screen[19][24] = 16'b10001_101010_11100;
end_screen[19][25] = 16'b10001_101010_11100;
end_screen[19][26] = 16'b10001_101010_11100;
end_screen[19][27] = 16'b10001_101010_11100;
end_screen[19][28] = 16'b10001_101010_11100;
end_screen[19][29] = 16'b10001_101010_11100;
end_screen[19][30] = 16'b10001_101010_11100;
end_screen[19][31] = 16'b10001_101010_11100;
end_screen[19][32] = 16'b10001_101010_11100;
end_screen[19][33] = 16'b10001_101010_11100;
end_screen[19][34] = 16'b10001_101010_11100;
end_screen[19][35] = 16'b10001_101010_11100;
end_screen[19][36] = 16'b10001_101010_11100;
end_screen[19][37] = 16'b10001_101010_11100;
end_screen[19][38] = 16'b10001_101010_11100;
end_screen[19][39] = 16'b10001_101010_11100;
end_screen[19][40] = 16'b10001_101010_11100;
end_screen[19][41] = 16'b10001_101010_11100;
end_screen[19][42] = 16'b10001_101010_11100;
end_screen[19][43] = 16'b10001_101010_11100;
end_screen[19][44] = 16'b10001_101010_11100;
end_screen[19][45] = 16'b10001_101010_11100;
end_screen[19][46] = 16'b10001_101010_11100;
end_screen[19][47] = 16'b10001_101010_11100;
end_screen[19][48] = 16'b10001_101010_11100;
end_screen[19][49] = 16'b10001_101010_11100;
end_screen[19][50] = 16'b10001_101010_11100;
end_screen[19][51] = 16'b10001_101010_11100;
end_screen[19][52] = 16'b10001_101010_11100;
end_screen[19][53] = 16'b10001_101010_11100;
end_screen[19][54] = 16'b10001_101010_11100;
end_screen[19][55] = 16'b10001_101010_11100;
end_screen[19][56] = 16'b10001_101010_11100;
end_screen[19][57] = 16'b10001_101010_11100;
end_screen[19][58] = 16'b10001_101010_11100;
end_screen[19][59] = 16'b10001_101010_11100;
end_screen[19][60] = 16'b10001_101010_11100;
end_screen[19][61] = 16'b10001_101010_11100;
end_screen[19][62] = 16'b10001_101010_11100;
end_screen[19][63] = 16'b10001_101010_11100;
end_screen[19][64] = 16'b10001_101010_11100;
end_screen[19][65] = 16'b10001_101010_11100;
end_screen[19][66] = 16'b10001_101010_11100;
end_screen[19][67] = 16'b10001_101010_11100;
end_screen[19][68] = 16'b10001_101010_11100;
end_screen[19][69] = 16'b10001_101010_11100;
end_screen[19][70] = 16'b10001_101010_11100;
end_screen[19][71] = 16'b10001_101010_11100;
end_screen[19][72] = 16'b10001_101010_11100;
end_screen[19][73] = 16'b10001_101010_11100;
end_screen[19][74] = 16'b10001_101010_11100;
end_screen[19][75] = 16'b10001_101010_11100;
end_screen[19][76] = 16'b10001_101010_11100;
end_screen[19][77] = 16'b10001_101010_11100;
end_screen[19][78] = 16'b10001_101010_11100;
end_screen[19][79] = 16'b10001_101010_11100;
end_screen[19][80] = 16'b10001_101010_11100;
end_screen[19][81] = 16'b10001_101010_11100;
end_screen[19][82] = 16'b10001_101010_11100;
end_screen[19][83] = 16'b10001_101010_11100;
end_screen[19][84] = 16'b10001_101010_11100;
end_screen[19][85] = 16'b10001_101010_11100;
end_screen[19][86] = 16'b10001_101010_11100;
end_screen[19][87] = 16'b10001_101010_11100;
end_screen[19][88] = 16'b10001_101010_11100;
end_screen[19][89] = 16'b10001_101010_11100;
end_screen[19][90] = 16'b10001_101010_11100;
end_screen[19][91] = 16'b10001_101010_11100;
end_screen[19][92] = 16'b10001_101010_11100;
end_screen[19][93] = 16'b10001_101010_11100;
end_screen[19][94] = 16'b10001_101010_11100;
end_screen[19][95] = 16'b10001_101010_11100;
end_screen[20][0] = 16'b10001_101010_11100;
end_screen[20][1] = 16'b10001_101010_11100;
end_screen[20][2] = 16'b10001_101010_11100;
end_screen[20][3] = 16'b10001_101010_11100;
end_screen[20][4] = 16'b10001_101010_11100;
end_screen[20][5] = 16'b10001_101010_11100;
end_screen[20][6] = 16'b10001_101010_11100;
end_screen[20][7] = 16'b10001_101010_11100;
end_screen[20][8] = 16'b10001_101010_11100;
end_screen[20][9] = 16'b10001_101010_11100;
end_screen[20][10] = 16'b10001_101010_11100;
end_screen[20][11] = 16'b10001_101010_11100;
end_screen[20][12] = 16'b10001_101010_11100;
end_screen[20][13] = 16'b10001_101010_11100;
end_screen[20][14] = 16'b10001_101010_11100;
end_screen[20][15] = 16'b10001_101010_11100;
end_screen[20][16] = 16'b10001_101010_11100;
end_screen[20][17] = 16'b10001_101010_11100;
end_screen[20][18] = 16'b10001_101010_11100;
end_screen[20][19] = 16'b10001_101010_11100;
end_screen[20][20] = 16'b10001_101010_11100;
end_screen[20][21] = 16'b10001_101010_11100;
end_screen[20][22] = 16'b10001_101010_11100;
end_screen[20][23] = 16'b10001_101010_11100;
end_screen[20][24] = 16'b10001_101010_11100;
end_screen[20][25] = 16'b10001_101010_11100;
end_screen[20][26] = 16'b10001_101010_11100;
end_screen[20][27] = 16'b10001_101010_11100;
end_screen[20][28] = 16'b10001_101010_11100;
end_screen[20][29] = 16'b10001_101010_11100;
end_screen[20][30] = 16'b10001_101010_11100;
end_screen[20][31] = 16'b10001_101010_11100;
end_screen[20][32] = 16'b10001_101010_11100;
end_screen[20][33] = 16'b10001_101010_11100;
end_screen[20][34] = 16'b10001_101010_11100;
end_screen[20][35] = 16'b10001_101010_11100;
end_screen[20][36] = 16'b10001_101010_11100;
end_screen[20][37] = 16'b10001_101010_11100;
end_screen[20][38] = 16'b10001_101010_11100;
end_screen[20][39] = 16'b10001_101010_11100;
end_screen[20][40] = 16'b10001_101010_11100;
end_screen[20][41] = 16'b10001_101010_11100;
end_screen[20][42] = 16'b10001_101010_11100;
end_screen[20][43] = 16'b10001_101010_11100;
end_screen[20][44] = 16'b10001_101010_11100;
end_screen[20][45] = 16'b10001_101010_11100;
end_screen[20][46] = 16'b10001_101010_11100;
end_screen[20][47] = 16'b10001_101010_11100;
end_screen[20][48] = 16'b10001_101010_11100;
end_screen[20][49] = 16'b10001_101010_11100;
end_screen[20][50] = 16'b10001_101010_11100;
end_screen[20][51] = 16'b10001_101010_11100;
end_screen[20][52] = 16'b10001_101010_11100;
end_screen[20][53] = 16'b10001_101010_11100;
end_screen[20][54] = 16'b10001_101010_11100;
end_screen[20][55] = 16'b10001_101010_11100;
end_screen[20][56] = 16'b10001_101010_11100;
end_screen[20][57] = 16'b10001_101010_11100;
end_screen[20][58] = 16'b10001_101010_11100;
end_screen[20][59] = 16'b10001_101010_11100;
end_screen[20][60] = 16'b10001_101010_11100;
end_screen[20][61] = 16'b10001_101010_11100;
end_screen[20][62] = 16'b10001_101010_11100;
end_screen[20][63] = 16'b10001_101010_11100;
end_screen[20][64] = 16'b10001_101010_11100;
end_screen[20][65] = 16'b10001_101010_11100;
end_screen[20][66] = 16'b10001_101010_11100;
end_screen[20][67] = 16'b10001_101010_11100;
end_screen[20][68] = 16'b10001_101010_11100;
end_screen[20][69] = 16'b10001_101010_11100;
end_screen[20][70] = 16'b10001_101010_11100;
end_screen[20][71] = 16'b10001_101010_11100;
end_screen[20][72] = 16'b10001_101010_11100;
end_screen[20][73] = 16'b10001_101010_11100;
end_screen[20][74] = 16'b10001_101010_11100;
end_screen[20][75] = 16'b10001_101010_11100;
end_screen[20][76] = 16'b10001_101010_11100;
end_screen[20][77] = 16'b10001_101010_11100;
end_screen[20][78] = 16'b10001_101010_11100;
end_screen[20][79] = 16'b10001_101010_11100;
end_screen[20][80] = 16'b10001_101010_11100;
end_screen[20][81] = 16'b10001_101010_11100;
end_screen[20][82] = 16'b10001_101010_11100;
end_screen[20][83] = 16'b10001_101010_11100;
end_screen[20][84] = 16'b10001_101010_11100;
end_screen[20][85] = 16'b10001_101010_11100;
end_screen[20][86] = 16'b10001_101010_11100;
end_screen[20][87] = 16'b10001_101010_11100;
end_screen[20][88] = 16'b10001_101010_11100;
end_screen[20][89] = 16'b10001_101010_11100;
end_screen[20][90] = 16'b10001_101010_11100;
end_screen[20][91] = 16'b10001_101010_11100;
end_screen[20][92] = 16'b10001_101010_11100;
end_screen[20][93] = 16'b10001_101010_11100;
end_screen[20][94] = 16'b10001_101010_11100;
end_screen[20][95] = 16'b10001_101010_11100;
end_screen[21][0] = 16'b10001_101010_11100;
end_screen[21][1] = 16'b10001_101010_11100;
end_screen[21][2] = 16'b10001_101010_11100;
end_screen[21][3] = 16'b10001_101010_11100;
end_screen[21][4] = 16'b10001_101010_11100;
end_screen[21][5] = 16'b10001_101010_11100;
end_screen[21][6] = 16'b10001_101010_11100;
end_screen[21][7] = 16'b10001_101010_11100;
end_screen[21][8] = 16'b10001_101010_11100;
end_screen[21][9] = 16'b10001_101010_11100;
end_screen[21][10] = 16'b10001_101010_11100;
end_screen[21][11] = 16'b10001_101010_11100;
end_screen[21][12] = 16'b10001_101010_11100;
end_screen[21][13] = 16'b10001_101010_11100;
end_screen[21][14] = 16'b10001_101010_11100;
end_screen[21][15] = 16'b10001_101010_11100;
end_screen[21][16] = 16'b10001_101010_11100;
end_screen[21][17] = 16'b10001_101010_11100;
end_screen[21][18] = 16'b10001_101010_11100;
end_screen[21][19] = 16'b10001_101010_11100;
end_screen[21][20] = 16'b10001_101010_11100;
end_screen[21][21] = 16'b10001_101010_11100;
end_screen[21][22] = 16'b10001_101010_11100;
end_screen[21][23] = 16'b10001_101010_11100;
end_screen[21][24] = 16'b10001_101010_11100;
end_screen[21][25] = 16'b10001_101010_11100;
end_screen[21][26] = 16'b10001_101010_11100;
end_screen[21][27] = 16'b10001_101010_11100;
end_screen[21][28] = 16'b10001_101010_11100;
end_screen[21][29] = 16'b10001_101010_11100;
end_screen[21][30] = 16'b10001_101010_11100;
end_screen[21][31] = 16'b10001_101010_11100;
end_screen[21][32] = 16'b10001_101010_11100;
end_screen[21][33] = 16'b10001_101010_11100;
end_screen[21][34] = 16'b10001_101010_11100;
end_screen[21][35] = 16'b10001_101010_11100;
end_screen[21][36] = 16'b10001_101010_11100;
end_screen[21][37] = 16'b10001_101010_11100;
end_screen[21][38] = 16'b10001_101010_11100;
end_screen[21][39] = 16'b10001_101010_11100;
end_screen[21][40] = 16'b10001_101010_11100;
end_screen[21][41] = 16'b10001_101010_11100;
end_screen[21][42] = 16'b10001_101010_11100;
end_screen[21][43] = 16'b10001_101010_11100;
end_screen[21][44] = 16'b10001_101010_11100;
end_screen[21][45] = 16'b10001_101010_11100;
end_screen[21][46] = 16'b10001_101010_11100;
end_screen[21][47] = 16'b10001_101010_11100;
end_screen[21][48] = 16'b10001_101010_11100;
end_screen[21][49] = 16'b10001_101010_11100;
end_screen[21][50] = 16'b10001_101010_11100;
end_screen[21][51] = 16'b10001_101010_11100;
end_screen[21][52] = 16'b10001_101010_11100;
end_screen[21][53] = 16'b10001_101010_11100;
end_screen[21][54] = 16'b10001_101010_11100;
end_screen[21][55] = 16'b10001_101010_11100;
end_screen[21][56] = 16'b10001_101010_11100;
end_screen[21][57] = 16'b10001_101010_11100;
end_screen[21][58] = 16'b10001_101010_11100;
end_screen[21][59] = 16'b10001_101010_11100;
end_screen[21][60] = 16'b10001_101010_11100;
end_screen[21][61] = 16'b10001_101010_11100;
end_screen[21][62] = 16'b10001_101010_11100;
end_screen[21][63] = 16'b10001_101010_11100;
end_screen[21][64] = 16'b10001_101010_11100;
end_screen[21][65] = 16'b10001_101010_11100;
end_screen[21][66] = 16'b10001_101010_11100;
end_screen[21][67] = 16'b10001_101010_11100;
end_screen[21][68] = 16'b10001_101010_11100;
end_screen[21][69] = 16'b10001_101010_11100;
end_screen[21][70] = 16'b10001_101010_11100;
end_screen[21][71] = 16'b10001_101010_11100;
end_screen[21][72] = 16'b10001_101010_11100;
end_screen[21][73] = 16'b10001_101010_11100;
end_screen[21][74] = 16'b10001_101010_11100;
end_screen[21][75] = 16'b10001_101010_11100;
end_screen[21][76] = 16'b10001_101010_11100;
end_screen[21][77] = 16'b10001_101010_11100;
end_screen[21][78] = 16'b10001_101010_11100;
end_screen[21][79] = 16'b10001_101010_11100;
end_screen[21][80] = 16'b10001_101010_11100;
end_screen[21][81] = 16'b10001_101010_11100;
end_screen[21][82] = 16'b10001_101010_11100;
end_screen[21][83] = 16'b10001_101010_11100;
end_screen[21][84] = 16'b10001_101010_11100;
end_screen[21][85] = 16'b10001_101010_11100;
end_screen[21][86] = 16'b10001_101010_11100;
end_screen[21][87] = 16'b10001_101010_11100;
end_screen[21][88] = 16'b10001_101010_11100;
end_screen[21][89] = 16'b10001_101010_11100;
end_screen[21][90] = 16'b10001_101010_11100;
end_screen[21][91] = 16'b10001_101010_11100;
end_screen[21][92] = 16'b10001_101010_11100;
end_screen[21][93] = 16'b10001_101010_11100;
end_screen[21][94] = 16'b10001_101010_11100;
end_screen[21][95] = 16'b10001_101010_11100;
end_screen[22][0] = 16'b10001_101010_11100;
end_screen[22][1] = 16'b10001_101010_11100;
end_screen[22][2] = 16'b10001_101010_11100;
end_screen[22][3] = 16'b10001_101010_11100;
end_screen[22][4] = 16'b10001_101010_11100;
end_screen[22][5] = 16'b10001_101010_11100;
end_screen[22][6] = 16'b10001_101010_11100;
end_screen[22][7] = 16'b10001_101010_11100;
end_screen[22][8] = 16'b10001_101010_11100;
end_screen[22][9] = 16'b10001_101010_11100;
end_screen[22][10] = 16'b10001_101010_11100;
end_screen[22][11] = 16'b10001_101010_11100;
end_screen[22][12] = 16'b10001_101010_11100;
end_screen[22][13] = 16'b10001_101010_11100;
end_screen[22][14] = 16'b10001_101010_11100;
end_screen[22][15] = 16'b10001_101010_11100;
end_screen[22][16] = 16'b10001_101010_11100;
end_screen[22][17] = 16'b10001_101010_11100;
end_screen[22][18] = 16'b10001_101010_11100;
end_screen[22][19] = 16'b10001_101010_11100;
end_screen[22][20] = 16'b10001_101010_11100;
end_screen[22][21] = 16'b10001_101010_11100;
end_screen[22][22] = 16'b10001_101010_11100;
end_screen[22][23] = 16'b10001_101010_11100;
end_screen[22][24] = 16'b10001_101010_11100;
end_screen[22][25] = 16'b10001_101010_11100;
end_screen[22][26] = 16'b10001_101010_11100;
end_screen[22][27] = 16'b10001_101010_11100;
end_screen[22][28] = 16'b10001_101010_11100;
end_screen[22][29] = 16'b10001_101010_11100;
end_screen[22][30] = 16'b10001_101010_11100;
end_screen[22][31] = 16'b10001_101010_11100;
end_screen[22][32] = 16'b10001_101010_11100;
end_screen[22][33] = 16'b10001_101010_11100;
end_screen[22][34] = 16'b10001_101010_11100;
end_screen[22][35] = 16'b10001_101010_11100;
end_screen[22][36] = 16'b10001_101010_11100;
end_screen[22][37] = 16'b10001_101010_11100;
end_screen[22][38] = 16'b10001_101010_11100;
end_screen[22][39] = 16'b10001_101010_11100;
end_screen[22][40] = 16'b10001_101010_11100;
end_screen[22][41] = 16'b10001_101010_11100;
end_screen[22][42] = 16'b10001_101010_11100;
end_screen[22][43] = 16'b10001_101010_11100;
end_screen[22][44] = 16'b10001_101010_11100;
end_screen[22][45] = 16'b10001_101010_11100;
end_screen[22][46] = 16'b10001_101010_11100;
end_screen[22][47] = 16'b10001_101010_11100;
end_screen[22][48] = 16'b10001_101010_11100;
end_screen[22][49] = 16'b10001_101010_11100;
end_screen[22][50] = 16'b10001_101010_11100;
end_screen[22][51] = 16'b10001_101010_11100;
end_screen[22][52] = 16'b10001_101010_11100;
end_screen[22][53] = 16'b10001_101010_11100;
end_screen[22][54] = 16'b10001_101010_11100;
end_screen[22][55] = 16'b10001_101010_11100;
end_screen[22][56] = 16'b10001_101010_11100;
end_screen[22][57] = 16'b10001_101010_11100;
end_screen[22][58] = 16'b10001_101010_11100;
end_screen[22][59] = 16'b10001_101010_11100;
end_screen[22][60] = 16'b10001_101010_11100;
end_screen[22][61] = 16'b10001_101010_11100;
end_screen[22][62] = 16'b10001_101010_11100;
end_screen[22][63] = 16'b10001_101010_11100;
end_screen[22][64] = 16'b10001_101010_11100;
end_screen[22][65] = 16'b10001_101010_11100;
end_screen[22][66] = 16'b10001_101010_11100;
end_screen[22][67] = 16'b10001_101010_11100;
end_screen[22][68] = 16'b10001_101010_11100;
end_screen[22][69] = 16'b10001_101010_11100;
end_screen[22][70] = 16'b10001_101010_11100;
end_screen[22][71] = 16'b10001_101010_11100;
end_screen[22][72] = 16'b10001_101010_11100;
end_screen[22][73] = 16'b10001_101010_11100;
end_screen[22][74] = 16'b10001_101010_11100;
end_screen[22][75] = 16'b10001_101010_11100;
end_screen[22][76] = 16'b10001_101010_11100;
end_screen[22][77] = 16'b10001_101010_11100;
end_screen[22][78] = 16'b10001_101010_11100;
end_screen[22][79] = 16'b10001_101010_11100;
end_screen[22][80] = 16'b10001_101010_11100;
end_screen[22][81] = 16'b10001_101010_11100;
end_screen[22][82] = 16'b10001_101010_11100;
end_screen[22][83] = 16'b10001_101010_11100;
end_screen[22][84] = 16'b10001_101010_11100;
end_screen[22][85] = 16'b10001_101010_11100;
end_screen[22][86] = 16'b10001_101010_11100;
end_screen[22][87] = 16'b10001_101010_11100;
end_screen[22][88] = 16'b10001_101010_11100;
end_screen[22][89] = 16'b10001_101010_11100;
end_screen[22][90] = 16'b10001_101010_11100;
end_screen[22][91] = 16'b10001_101010_11100;
end_screen[22][92] = 16'b10001_101010_11100;
end_screen[22][93] = 16'b10001_101010_11100;
end_screen[22][94] = 16'b10001_101010_11100;
end_screen[22][95] = 16'b10001_101010_11100;
end_screen[23][0] = 16'b10001_101010_11100;
end_screen[23][1] = 16'b10001_101010_11100;
end_screen[23][2] = 16'b10001_101010_11100;
end_screen[23][3] = 16'b10001_101010_11100;
end_screen[23][4] = 16'b10001_101010_11100;
end_screen[23][5] = 16'b10001_101010_11100;
end_screen[23][6] = 16'b10001_101010_11100;
end_screen[23][7] = 16'b10001_101010_11100;
end_screen[23][8] = 16'b10001_101010_11100;
end_screen[23][9] = 16'b10001_101010_11100;
end_screen[23][10] = 16'b10001_101010_11100;
end_screen[23][11] = 16'b10001_101010_11100;
end_screen[23][12] = 16'b10001_101010_11100;
end_screen[23][13] = 16'b10001_101010_11100;
end_screen[23][14] = 16'b10001_101010_11100;
end_screen[23][15] = 16'b10001_101010_11100;
end_screen[23][16] = 16'b10001_101010_11100;
end_screen[23][17] = 16'b10001_101010_11100;
end_screen[23][18] = 16'b10001_101010_11100;
end_screen[23][19] = 16'b10001_101010_11100;
end_screen[23][20] = 16'b10001_101010_11100;
end_screen[23][21] = 16'b10001_101010_11100;
end_screen[23][22] = 16'b10001_101010_11100;
end_screen[23][23] = 16'b10001_101010_11100;
end_screen[23][24] = 16'b10001_101010_11100;
end_screen[23][25] = 16'b10001_101010_11100;
end_screen[23][26] = 16'b10001_101010_11100;
end_screen[23][27] = 16'b10001_101010_11100;
end_screen[23][28] = 16'b10001_101010_11100;
end_screen[23][29] = 16'b10001_101010_11100;
end_screen[23][30] = 16'b10001_101010_11100;
end_screen[23][31] = 16'b10001_101010_11100;
end_screen[23][32] = 16'b10010_101010_11011;
end_screen[23][33] = 16'b10010_101010_11011;
end_screen[23][34] = 16'b10010_101010_11011;
end_screen[23][35] = 16'b10001_101001_11011;
end_screen[23][36] = 16'b10010_101010_11011;
end_screen[23][37] = 16'b10010_101010_11011;
end_screen[23][38] = 16'b10010_101010_11011;
end_screen[23][39] = 16'b10010_101010_11011;
end_screen[23][40] = 16'b10010_101010_11011;
end_screen[23][41] = 16'b10010_101010_11011;
end_screen[23][42] = 16'b10010_101010_11011;
end_screen[23][43] = 16'b10010_101010_11011;
end_screen[23][44] = 16'b10010_101010_11011;
end_screen[23][45] = 16'b10010_101011_11011;
end_screen[23][46] = 16'b10001_101010_11100;
end_screen[23][47] = 16'b10001_101010_11100;
end_screen[23][48] = 16'b10001_101010_11100;
end_screen[23][49] = 16'b10001_101010_11100;
end_screen[23][50] = 16'b10001_101010_11100;
end_screen[23][51] = 16'b10001_101010_11100;
end_screen[23][52] = 16'b10001_101010_11100;
end_screen[23][53] = 16'b10001_101010_11100;
end_screen[23][54] = 16'b10001_101010_11100;
end_screen[23][55] = 16'b10001_101010_11100;
end_screen[23][56] = 16'b10001_101010_11100;
end_screen[23][57] = 16'b10001_101010_11100;
end_screen[23][58] = 16'b10001_101010_11100;
end_screen[23][59] = 16'b10101_100101_10100;
end_screen[23][60] = 16'b10111_011111_01101;
end_screen[23][61] = 16'b10111_011111_01110;
end_screen[23][62] = 16'b10111_100000_01110;
end_screen[23][63] = 16'b10111_011111_01110;
end_screen[23][64] = 16'b10111_011111_01110;
end_screen[23][65] = 16'b10101_100010_10011;
end_screen[23][66] = 16'b10001_101010_11100;
end_screen[23][67] = 16'b10001_101010_11100;
end_screen[23][68] = 16'b10001_101010_11100;
end_screen[23][69] = 16'b10001_101010_11100;
end_screen[23][70] = 16'b10001_101010_11100;
end_screen[23][71] = 16'b10001_101010_11100;
end_screen[23][72] = 16'b10001_101010_11100;
end_screen[23][73] = 16'b10001_101010_11100;
end_screen[23][74] = 16'b10001_101010_11100;
end_screen[23][75] = 16'b10001_101010_11100;
end_screen[23][76] = 16'b10001_101010_11100;
end_screen[23][77] = 16'b10001_101010_11100;
end_screen[23][78] = 16'b10001_101010_11100;
end_screen[23][79] = 16'b10001_101010_11100;
end_screen[23][80] = 16'b10001_101010_11100;
end_screen[23][81] = 16'b10001_101010_11100;
end_screen[23][82] = 16'b10001_101010_11100;
end_screen[23][83] = 16'b10001_101010_11100;
end_screen[23][84] = 16'b10001_101010_11100;
end_screen[23][85] = 16'b10001_101010_11100;
end_screen[23][86] = 16'b10001_101010_11100;
end_screen[23][87] = 16'b10001_101010_11100;
end_screen[23][88] = 16'b10001_101010_11100;
end_screen[23][89] = 16'b10001_101010_11100;
end_screen[23][90] = 16'b10001_101010_11100;
end_screen[23][91] = 16'b10001_101010_11100;
end_screen[23][92] = 16'b10001_101010_11100;
end_screen[23][93] = 16'b10001_101010_11100;
end_screen[23][94] = 16'b10001_101010_11100;
end_screen[23][95] = 16'b10001_101010_11100;
end_screen[24][0] = 16'b10001_101010_11100;
end_screen[24][1] = 16'b10001_101010_11100;
end_screen[24][2] = 16'b10001_101010_11100;
end_screen[24][3] = 16'b10001_101010_11100;
end_screen[24][4] = 16'b10001_101010_11100;
end_screen[24][5] = 16'b10001_101010_11100;
end_screen[24][6] = 16'b10001_101010_11100;
end_screen[24][7] = 16'b10001_101010_11100;
end_screen[24][8] = 16'b10001_101010_11100;
end_screen[24][9] = 16'b10001_101010_11100;
end_screen[24][10] = 16'b10001_101010_11100;
end_screen[24][11] = 16'b10001_101010_11100;
end_screen[24][12] = 16'b10001_101010_11100;
end_screen[24][13] = 16'b10001_101010_11100;
end_screen[24][14] = 16'b10001_101010_11100;
end_screen[24][15] = 16'b10001_101010_11100;
end_screen[24][16] = 16'b10001_101010_11100;
end_screen[24][17] = 16'b10001_101010_11100;
end_screen[24][18] = 16'b10001_101010_11100;
end_screen[24][19] = 16'b10001_101010_11100;
end_screen[24][20] = 16'b10001_101010_11100;
end_screen[24][21] = 16'b10001_101010_11100;
end_screen[24][22] = 16'b10001_101010_11100;
end_screen[24][23] = 16'b10001_101010_11100;
end_screen[24][24] = 16'b10001_101010_11100;
end_screen[24][25] = 16'b10001_101010_11100;
end_screen[24][26] = 16'b10001_101010_11100;
end_screen[24][27] = 16'b10001_101010_11100;
end_screen[24][28] = 16'b10001_101010_11100;
end_screen[24][29] = 16'b10001_101010_11100;
end_screen[24][30] = 16'b10001_101010_11100;
end_screen[24][31] = 16'b10101_101001_10101;
end_screen[24][32] = 16'b11010_101010_01110;
end_screen[24][33] = 16'b11000_100100_01011;
end_screen[24][34] = 16'b10001_010101_00011;
end_screen[24][35] = 16'b10001_010101_00011;
end_screen[24][36] = 16'b10011_011000_00101;
end_screen[24][37] = 16'b10100_011010_00101;
end_screen[24][38] = 16'b10100_011011_00110;
end_screen[24][39] = 16'b10100_011011_00110;
end_screen[24][40] = 16'b10100_011011_00110;
end_screen[24][41] = 16'b10100_011010_00101;
end_screen[24][42] = 16'b10011_011001_00101;
end_screen[24][43] = 16'b10011_010111_00100;
end_screen[24][44] = 16'b11000_100100_01011;
end_screen[24][45] = 16'b11010_101011_01110;
end_screen[24][46] = 16'b10101_101010_10101;
end_screen[24][47] = 16'b10001_101010_11100;
end_screen[24][48] = 16'b10001_101010_11100;
end_screen[24][49] = 16'b10001_101010_11100;
end_screen[24][50] = 16'b10001_101010_11100;
end_screen[24][51] = 16'b10001_101010_11100;
end_screen[24][52] = 16'b10001_101010_11100;
end_screen[24][53] = 16'b10001_101010_11100;
end_screen[24][54] = 16'b10001_101010_11100;
end_screen[24][55] = 16'b10001_101010_11100;
end_screen[24][56] = 16'b10001_101010_11100;
end_screen[24][57] = 16'b10101_101000_10101;
end_screen[24][58] = 16'b10110_100110_10011;
end_screen[24][59] = 16'b11011_011010_00101;
end_screen[24][60] = 16'b11100_010111_00011;
end_screen[24][61] = 16'b11100_011000_00011;
end_screen[24][62] = 16'b11100_011000_00011;
end_screen[24][63] = 16'b11100_011000_00011;
end_screen[24][64] = 16'b11100_010111_00011;
end_screen[24][65] = 16'b11011_011000_00100;
end_screen[24][66] = 16'b10110_100100_10010;
end_screen[24][67] = 16'b10101_100011_10010;
end_screen[24][68] = 16'b10001_101010_11100;
end_screen[24][69] = 16'b10001_101010_11100;
end_screen[24][70] = 16'b10001_101010_11100;
end_screen[24][71] = 16'b10001_101010_11100;
end_screen[24][72] = 16'b10001_101010_11100;
end_screen[24][73] = 16'b10001_101010_11100;
end_screen[24][74] = 16'b10001_101010_11100;
end_screen[24][75] = 16'b10001_101010_11100;
end_screen[24][76] = 16'b10001_101010_11100;
end_screen[24][77] = 16'b10001_101010_11100;
end_screen[24][78] = 16'b10001_101010_11100;
end_screen[24][79] = 16'b10001_101010_11100;
end_screen[24][80] = 16'b10001_101010_11100;
end_screen[24][81] = 16'b10001_101010_11100;
end_screen[24][82] = 16'b10001_101010_11100;
end_screen[24][83] = 16'b10001_101010_11100;
end_screen[24][84] = 16'b10001_101010_11100;
end_screen[24][85] = 16'b10001_101010_11100;
end_screen[24][86] = 16'b10001_101010_11100;
end_screen[24][87] = 16'b10001_101010_11100;
end_screen[24][88] = 16'b10001_101010_11100;
end_screen[24][89] = 16'b10001_101010_11100;
end_screen[24][90] = 16'b10001_101010_11100;
end_screen[24][91] = 16'b10001_101010_11100;
end_screen[24][92] = 16'b10001_101010_11100;
end_screen[24][93] = 16'b10001_101010_11100;
end_screen[24][94] = 16'b10001_101010_11100;
end_screen[24][95] = 16'b10001_101010_11100;
end_screen[25][0] = 16'b10001_101010_11100;
end_screen[25][1] = 16'b10001_101010_11100;
end_screen[25][2] = 16'b10001_101010_11100;
end_screen[25][3] = 16'b10001_101010_11100;
end_screen[25][4] = 16'b10001_101010_11100;
end_screen[25][5] = 16'b10001_101010_11100;
end_screen[25][6] = 16'b10001_101010_11100;
end_screen[25][7] = 16'b10001_101010_11100;
end_screen[25][8] = 16'b10001_101010_11100;
end_screen[25][9] = 16'b10001_101010_11100;
end_screen[25][10] = 16'b10001_101010_11100;
end_screen[25][11] = 16'b10001_101010_11100;
end_screen[25][12] = 16'b10001_101010_11100;
end_screen[25][13] = 16'b10001_101010_11100;
end_screen[25][14] = 16'b10001_101010_11100;
end_screen[25][15] = 16'b10001_101010_11100;
end_screen[25][16] = 16'b10001_101010_11100;
end_screen[25][17] = 16'b10001_101010_11100;
end_screen[25][18] = 16'b10001_101010_11100;
end_screen[25][19] = 16'b10001_101010_11100;
end_screen[25][20] = 16'b10001_101010_11100;
end_screen[25][21] = 16'b10001_101010_11100;
end_screen[25][22] = 16'b10001_101010_11100;
end_screen[25][23] = 16'b10001_101010_11100;
end_screen[25][24] = 16'b10001_101010_11100;
end_screen[25][25] = 16'b10001_101010_11100;
end_screen[25][26] = 16'b10001_101010_11100;
end_screen[25][27] = 16'b10001_101010_11100;
end_screen[25][28] = 16'b10001_101010_11100;
end_screen[25][29] = 16'b10100_100011_01110;
end_screen[25][30] = 16'b10010_011010_00110;
end_screen[25][31] = 16'b10010_010111_00100;
end_screen[25][32] = 16'b10100_011010_00101;
end_screen[25][33] = 16'b10101_011100_00101;
end_screen[25][34] = 16'b10110_011101_00110;
end_screen[25][35] = 16'b10101_011101_00110;
end_screen[25][36] = 16'b10110_011101_00110;
end_screen[25][37] = 16'b10110_011110_00110;
end_screen[25][38] = 16'b10110_011110_00110;
end_screen[25][39] = 16'b10111_011111_00111;
end_screen[25][40] = 16'b10111_100000_00111;
end_screen[25][41] = 16'b10111_100000_00111;
end_screen[25][42] = 16'b10110_011110_00110;
end_screen[25][43] = 16'b10101_011100_00101;
end_screen[25][44] = 16'b10101_011011_00101;
end_screen[25][45] = 16'b10011_011001_00100;
end_screen[25][46] = 16'b10011_011000_00100;
end_screen[25][47] = 16'b10100_011100_00111;
end_screen[25][48] = 16'b10101_100110_10001;
end_screen[25][49] = 16'b10001_101010_11100;
end_screen[25][50] = 16'b10001_101010_11100;
end_screen[25][51] = 16'b10001_101010_11100;
end_screen[25][52] = 16'b10001_101010_11100;
end_screen[25][53] = 16'b10001_101010_11100;
end_screen[25][54] = 16'b10001_101010_11100;
end_screen[25][55] = 16'b10001_101010_11100;
end_screen[25][56] = 16'b10101_100100_10011;
end_screen[25][57] = 16'b11100_011100_00110;
end_screen[25][58] = 16'b11100_011011_00100;
end_screen[25][59] = 16'b11100_011001_00100;
end_screen[25][60] = 16'b11011_011000_00100;
end_screen[25][61] = 16'b11011_010111_00011;
end_screen[25][62] = 16'b11011_010111_00011;
end_screen[25][63] = 16'b11100_011010_00100;
end_screen[25][64] = 16'b11100_011010_00100;
end_screen[25][65] = 16'b11100_011011_00101;
end_screen[25][66] = 16'b11011_010110_00010;
end_screen[25][67] = 16'b11011_010010_00001;
end_screen[25][68] = 16'b10110_100000_10000;
end_screen[25][69] = 16'b10110_100110_10011;
end_screen[25][70] = 16'b10010_101001_11011;
end_screen[25][71] = 16'b10001_101010_11100;
end_screen[25][72] = 16'b10001_101010_11100;
end_screen[25][73] = 16'b10001_101010_11100;
end_screen[25][74] = 16'b10001_101010_11100;
end_screen[25][75] = 16'b10001_101010_11100;
end_screen[25][76] = 16'b10001_101010_11100;
end_screen[25][77] = 16'b10001_101010_11100;
end_screen[25][78] = 16'b10001_101010_11100;
end_screen[25][79] = 16'b10001_101010_11100;
end_screen[25][80] = 16'b10001_101010_11100;
end_screen[25][81] = 16'b10001_101010_11100;
end_screen[25][82] = 16'b10001_101010_11100;
end_screen[25][83] = 16'b10001_101010_11100;
end_screen[25][84] = 16'b10001_101010_11100;
end_screen[25][85] = 16'b10001_101010_11100;
end_screen[25][86] = 16'b10001_101010_11100;
end_screen[25][87] = 16'b10001_101010_11100;
end_screen[25][88] = 16'b10001_101010_11100;
end_screen[25][89] = 16'b10001_101010_11100;
end_screen[25][90] = 16'b10001_101010_11100;
end_screen[25][91] = 16'b10001_101010_11100;
end_screen[25][92] = 16'b10001_101010_11100;
end_screen[25][93] = 16'b10001_101010_11100;
end_screen[25][94] = 16'b10001_101010_11100;
end_screen[25][95] = 16'b10001_101010_11100;
end_screen[26][0] = 16'b10001_101010_11100;
end_screen[26][1] = 16'b10001_101010_11100;
end_screen[26][2] = 16'b10001_101010_11100;
end_screen[26][3] = 16'b10001_101010_11100;
end_screen[26][4] = 16'b10001_101010_11100;
end_screen[26][5] = 16'b10001_101010_11100;
end_screen[26][6] = 16'b10001_101010_11100;
end_screen[26][7] = 16'b10001_101010_11100;
end_screen[26][8] = 16'b10001_101010_11100;
end_screen[26][9] = 16'b10001_101010_11100;
end_screen[26][10] = 16'b10001_101010_11100;
end_screen[26][11] = 16'b10001_101010_11100;
end_screen[26][12] = 16'b10001_101010_11100;
end_screen[26][13] = 16'b10001_101010_11100;
end_screen[26][14] = 16'b10001_101010_11100;
end_screen[26][15] = 16'b10001_101010_11100;
end_screen[26][16] = 16'b10001_101010_11100;
end_screen[26][17] = 16'b10001_101010_11100;
end_screen[26][18] = 16'b10001_101010_11100;
end_screen[26][19] = 16'b10001_101010_11100;
end_screen[26][20] = 16'b10001_101010_11100;
end_screen[26][21] = 16'b10001_101010_11100;
end_screen[26][22] = 16'b10001_101010_11100;
end_screen[26][23] = 16'b10001_101010_11100;
end_screen[26][24] = 16'b10001_101010_11100;
end_screen[26][25] = 16'b10001_101010_11100;
end_screen[26][26] = 16'b10001_101010_11100;
end_screen[26][27] = 16'b10110_100100_01101;
end_screen[26][28] = 16'b10010_011100_01001;
end_screen[26][29] = 16'b10001_010100_00010;
end_screen[26][30] = 16'b10001_010100_00010;
end_screen[26][31] = 16'b10011_010111_00011;
end_screen[26][32] = 16'b10100_011001_00100;
end_screen[26][33] = 16'b10100_011010_00101;
end_screen[26][34] = 16'b10110_011111_00111;
end_screen[26][35] = 16'b10110_011110_00110;
end_screen[26][36] = 16'b10100_011011_00101;
end_screen[26][37] = 16'b10100_011011_00101;
end_screen[26][38] = 16'b11111_111111_11111;
end_screen[26][39] = 16'b11111_111111_11111;
end_screen[26][40] = 16'b11111_111111_11111;
end_screen[26][41] = 16'b11111_111111_11111;
end_screen[26][42] = 16'b11111_111111_11111;
end_screen[26][43] = 16'b11111_111111_11111;
end_screen[26][44] = 16'b11111_111111_11111;
end_screen[26][45] = 16'b11111_111111_11111;
end_screen[26][46] = 16'b11111_111111_11111;
end_screen[26][47] = 16'b11111_111111_11111;
end_screen[26][48] = 16'b11111_111111_11111;
end_screen[26][49] = 16'b11111_111111_11111;
end_screen[26][50] = 16'b11111_111111_11111;
end_screen[26][51] = 16'b11111_111111_11111;
end_screen[26][52] = 16'b11111_111111_11111;
end_screen[26][53] = 16'b11111_111111_11111;
end_screen[26][54] = 16'b11111_111111_11111;
end_screen[26][55] = 16'b11111_111111_11111;
end_screen[26][56] = 16'b11111_111111_11111;
end_screen[26][57] = 16'b11111_111111_11111;
end_screen[26][58] = 16'b11111_111111_11111;
end_screen[26][59] = 16'b11100_011010_00100;
end_screen[26][60] = 16'b11011_010110_00011;
end_screen[26][61] = 16'b11011_011000_00100;
end_screen[26][62] = 16'b11100_011011_00101;
end_screen[26][63] = 16'b11100_011001_00100;
end_screen[26][64] = 16'b11100_011001_00100;
end_screen[26][65] = 16'b11100_011101_00110;
end_screen[26][66] = 16'b11011_010111_00011;
end_screen[26][67] = 16'b11011_010100_00010;
end_screen[26][68] = 16'b11011_010110_00011;
end_screen[26][69] = 16'b11101_011101_00110;
end_screen[26][70] = 16'b10011_101000_11001;
end_screen[26][71] = 16'b10001_101010_11100;
end_screen[26][72] = 16'b10001_101010_11100;
end_screen[26][73] = 16'b10001_101010_11100;
end_screen[26][74] = 16'b10001_101010_11100;
end_screen[26][75] = 16'b10001_101010_11100;
end_screen[26][76] = 16'b10001_101010_11100;
end_screen[26][77] = 16'b10001_101010_11100;
end_screen[26][78] = 16'b10001_101010_11100;
end_screen[26][79] = 16'b10001_101010_11100;
end_screen[26][80] = 16'b10001_101010_11100;
end_screen[26][81] = 16'b10001_101010_11100;
end_screen[26][82] = 16'b10001_101010_11100;
end_screen[26][83] = 16'b10001_101010_11100;
end_screen[26][84] = 16'b10001_101010_11100;
end_screen[26][85] = 16'b10001_101010_11100;
end_screen[26][86] = 16'b10001_101010_11100;
end_screen[26][87] = 16'b10001_101010_11100;
end_screen[26][88] = 16'b10001_101010_11100;
end_screen[26][89] = 16'b10001_101010_11100;
end_screen[26][90] = 16'b10001_101010_11100;
end_screen[26][91] = 16'b10001_101010_11100;
end_screen[26][92] = 16'b10001_101010_11100;
end_screen[26][93] = 16'b10001_101010_11100;
end_screen[26][94] = 16'b10001_101010_11100;
end_screen[26][95] = 16'b10001_101010_11100;
end_screen[27][0] = 16'b10001_101010_11100;
end_screen[27][1] = 16'b10001_101010_11100;
end_screen[27][2] = 16'b10001_101010_11100;
end_screen[27][3] = 16'b10001_101010_11100;
end_screen[27][4] = 16'b10001_101010_11100;
end_screen[27][5] = 16'b10001_101010_11100;
end_screen[27][6] = 16'b10001_101010_11100;
end_screen[27][7] = 16'b10001_101010_11100;
end_screen[27][8] = 16'b10001_101010_11100;
end_screen[27][9] = 16'b10001_101010_11100;
end_screen[27][10] = 16'b10001_101010_11100;
end_screen[27][11] = 16'b10001_101010_11100;
end_screen[27][12] = 16'b10001_101010_11100;
end_screen[27][13] = 16'b10001_101010_11100;
end_screen[27][14] = 16'b10001_101010_11100;
end_screen[27][15] = 16'b10001_101010_11100;
end_screen[27][16] = 16'b10001_101010_11100;
end_screen[27][17] = 16'b10001_101010_11100;
end_screen[27][18] = 16'b10001_101010_11100;
end_screen[27][19] = 16'b10001_101010_11100;
end_screen[27][20] = 16'b10001_101010_11100;
end_screen[27][21] = 16'b10001_101010_11100;
end_screen[27][22] = 16'b10001_101010_11100;
end_screen[27][23] = 16'b10001_101010_11100;
end_screen[27][24] = 16'b10001_101010_11100;
end_screen[27][25] = 16'b10010_101001_11001;
end_screen[27][26] = 16'b10101_100010_01101;
end_screen[27][27] = 16'b10100_011010_00100;
end_screen[27][28] = 16'b10010_010110_00011;
end_screen[27][29] = 16'b10010_010110_00011;
end_screen[27][30] = 16'b10010_010111_00100;
end_screen[27][31] = 16'b10011_011000_00100;
end_screen[27][32] = 16'b10010_010110_00011;
end_screen[27][33] = 16'b10000_010011_00010;
end_screen[27][34] = 16'b01110_001111_00001;
end_screen[27][35] = 16'b01101_001110_00001;
end_screen[27][36] = 16'b01110_001111_00001;
end_screen[27][37] = 16'b01101_001110_00001;
end_screen[27][38] = 16'b11111_111111_11111;
end_screen[27][39] = 16'b11111_111111_11111;
end_screen[27][40] = 16'b11111_111111_11111;
end_screen[27][41] = 16'b11111_111111_11111;
end_screen[27][42] = 16'b11111_111111_11111;
end_screen[27][43] = 16'b11111_111111_11111;
end_screen[27][44] = 16'b11111_111111_11111;
end_screen[27][45] = 16'b11111_111111_11111;
end_screen[27][46] = 16'b11111_111111_11111;
end_screen[27][47] = 16'b11111_111111_11111;
end_screen[27][48] = 16'b11111_111111_11111;
end_screen[27][49] = 16'b11111_111111_11111;
end_screen[27][50] = 16'b11111_111111_11111;
end_screen[27][51] = 16'b11111_111111_11111;
end_screen[27][52] = 16'b11111_111111_11111;
end_screen[27][53] = 16'b11111_111111_11111;
end_screen[27][54] = 16'b11111_111111_11111;
end_screen[27][55] = 16'b11111_111111_11111;
end_screen[27][56] = 16'b11111_111111_11111;
end_screen[27][57] = 16'b11111_111111_11111;
end_screen[27][58] = 16'b11111_111111_11111;
end_screen[27][59] = 16'b11011_010110_00011;
end_screen[27][60] = 16'b11011_010100_00010;
end_screen[27][61] = 16'b11100_011001_00100;
end_screen[27][62] = 16'b11100_011110_00110;
end_screen[27][63] = 16'b11100_011011_00101;
end_screen[27][64] = 16'b11011_010101_00010;
end_screen[27][65] = 16'b11011_011000_00011;
end_screen[27][66] = 16'b11100_011001_00100;
end_screen[27][67] = 16'b11100_011011_00101;
end_screen[27][68] = 16'b11100_011001_00100;
end_screen[27][69] = 16'b11011_010100_00010;
end_screen[27][70] = 16'b10110_100001_01111;
end_screen[27][71] = 16'b10001_101010_11100;
end_screen[27][72] = 16'b10001_101010_11100;
end_screen[27][73] = 16'b10001_101010_11100;
end_screen[27][74] = 16'b10001_101010_11100;
end_screen[27][75] = 16'b10001_101010_11100;
end_screen[27][76] = 16'b10001_101010_11100;
end_screen[27][77] = 16'b10001_101010_11100;
end_screen[27][78] = 16'b10001_101010_11100;
end_screen[27][79] = 16'b10001_101010_11100;
end_screen[27][80] = 16'b10001_101010_11100;
end_screen[27][81] = 16'b10001_101010_11100;
end_screen[27][82] = 16'b10001_101010_11100;
end_screen[27][83] = 16'b10001_101010_11100;
end_screen[27][84] = 16'b10001_101010_11100;
end_screen[27][85] = 16'b10001_101010_11100;
end_screen[27][86] = 16'b10001_101010_11100;
end_screen[27][87] = 16'b10001_101010_11100;
end_screen[27][88] = 16'b10001_101010_11100;
end_screen[27][89] = 16'b10001_101010_11100;
end_screen[27][90] = 16'b10001_101010_11100;
end_screen[27][91] = 16'b10001_101010_11100;
end_screen[27][92] = 16'b10001_101010_11100;
end_screen[27][93] = 16'b10001_101010_11100;
end_screen[27][94] = 16'b10001_101010_11100;
end_screen[27][95] = 16'b10001_101010_11100;
end_screen[28][0] = 16'b10001_101010_11100;
end_screen[28][1] = 16'b10001_101010_11100;
end_screen[28][2] = 16'b10001_101010_11100;
end_screen[28][3] = 16'b10001_101010_11100;
end_screen[28][4] = 16'b10001_101010_11100;
end_screen[28][5] = 16'b10001_101010_11100;
end_screen[28][6] = 16'b10001_101010_11100;
end_screen[28][7] = 16'b10001_101010_11100;
end_screen[28][8] = 16'b10001_101010_11100;
end_screen[28][9] = 16'b10001_101010_11100;
end_screen[28][10] = 16'b10001_101010_11100;
end_screen[28][11] = 16'b10001_101010_11100;
end_screen[28][12] = 16'b10001_101010_11100;
end_screen[28][13] = 16'b10001_101010_11100;
end_screen[28][14] = 16'b10001_101010_11100;
end_screen[28][15] = 16'b10001_101010_11100;
end_screen[28][16] = 16'b10001_101010_11100;
end_screen[28][17] = 16'b10001_101010_11100;
end_screen[28][18] = 16'b10001_101010_11100;
end_screen[28][19] = 16'b10001_101010_11100;
end_screen[28][20] = 16'b10001_101010_11100;
end_screen[28][21] = 16'b10001_101010_11100;
end_screen[28][22] = 16'b10001_101010_11100;
end_screen[28][23] = 16'b10001_101010_11100;
end_screen[28][24] = 16'b10001_101010_11100;
end_screen[28][25] = 16'b10010_101001_11001;
end_screen[28][26] = 16'b10010_010111_00011;
end_screen[28][27] = 16'b10011_010111_00100;
end_screen[28][28] = 16'b10100_011010_00101;
end_screen[28][29] = 16'b10000_010100_00011;
end_screen[28][30] = 16'b01110_010000_00010;
end_screen[28][31] = 16'b01110_010001_00010;
end_screen[28][32] = 16'b01110_001111_00001;
end_screen[28][33] = 16'b01011_001010_00000;
end_screen[28][34] = 16'b01001_001000_00000;
end_screen[28][35] = 16'b01010_001001_00001;
end_screen[28][36] = 16'b01100_001100_00001;
end_screen[28][37] = 16'b01010_001011_00001;
end_screen[28][38] = 16'b11111_111111_11111;
end_screen[28][39] = 16'b11111_111111_11111;
end_screen[28][40] = 16'b11111_111111_11111;
end_screen[28][41] = 16'b11111_111111_11111;
end_screen[28][42] = 16'b11111_111111_11111;
end_screen[28][43] = 16'b11111_111111_11111;
end_screen[28][44] = 16'b11111_111111_11111;
end_screen[28][45] = 16'b11111_111111_11111;
end_screen[28][46] = 16'b11111_111111_11111;
end_screen[28][47] = 16'b11111_111111_11111;
end_screen[28][48] = 16'b11111_111111_11111;
end_screen[28][49] = 16'b11111_111111_11111;
end_screen[28][50] = 16'b11111_111111_11111;
end_screen[28][51] = 16'b11111_111111_11111;
end_screen[28][52] = 16'b11111_111111_11111;
end_screen[28][53] = 16'b11111_111111_11111;
end_screen[28][54] = 16'b11111_111111_11111;
end_screen[28][55] = 16'b11111_111111_11111;
end_screen[28][56] = 16'b11111_111111_11111;
end_screen[28][57] = 16'b11111_111111_11111;
end_screen[28][58] = 16'b11111_111111_11111;
end_screen[28][59] = 16'b11011_011001_00100;
end_screen[28][60] = 16'b11100_011010_00100;
end_screen[28][61] = 16'b11011_010111_00011;
end_screen[28][62] = 16'b11100_011010_00100;
end_screen[28][63] = 16'b11100_011011_00101;
end_screen[28][64] = 16'b11011_010111_00011;
end_screen[28][65] = 16'b11011_010111_00011;
end_screen[28][66] = 16'b11100_011100_00101;
end_screen[28][67] = 16'b11011_011001_00100;
end_screen[28][68] = 16'b11011_010100_00010;
end_screen[28][69] = 16'b11010_010001_00001;
end_screen[28][70] = 16'b11011_010010_00001;
end_screen[28][71] = 16'b10111_100010_10000;
end_screen[28][72] = 16'b10001_101010_11100;
end_screen[28][73] = 16'b10001_101010_11100;
end_screen[28][74] = 16'b10001_101010_11100;
end_screen[28][75] = 16'b10001_101010_11100;
end_screen[28][76] = 16'b10001_101010_11100;
end_screen[28][77] = 16'b10001_101010_11100;
end_screen[28][78] = 16'b10001_101010_11100;
end_screen[28][79] = 16'b10001_101010_11100;
end_screen[28][80] = 16'b10001_101010_11100;
end_screen[28][81] = 16'b10001_101010_11100;
end_screen[28][82] = 16'b10001_101010_11100;
end_screen[28][83] = 16'b10001_101010_11100;
end_screen[28][84] = 16'b10001_101010_11100;
end_screen[28][85] = 16'b10001_101010_11100;
end_screen[28][86] = 16'b10001_101010_11100;
end_screen[28][87] = 16'b10001_101010_11100;
end_screen[28][88] = 16'b10001_101010_11100;
end_screen[28][89] = 16'b10001_101010_11100;
end_screen[28][90] = 16'b10001_101010_11100;
end_screen[28][91] = 16'b10001_101010_11100;
end_screen[28][92] = 16'b10001_101010_11100;
end_screen[28][93] = 16'b10001_101010_11100;
end_screen[28][94] = 16'b10001_101010_11100;
end_screen[28][95] = 16'b10001_101010_11100;
end_screen[29][0] = 16'b10001_101010_11100;
end_screen[29][1] = 16'b10001_101010_11100;
end_screen[29][2] = 16'b10001_101010_11100;
end_screen[29][3] = 16'b10001_101010_11100;
end_screen[29][4] = 16'b10001_101010_11100;
end_screen[29][5] = 16'b10001_101010_11100;
end_screen[29][6] = 16'b10001_101010_11100;
end_screen[29][7] = 16'b10001_101010_11100;
end_screen[29][8] = 16'b10001_101010_11100;
end_screen[29][9] = 16'b10001_101010_11100;
end_screen[29][10] = 16'b10001_101010_11100;
end_screen[29][11] = 16'b10001_101010_11100;
end_screen[29][12] = 16'b10001_101010_11100;
end_screen[29][13] = 16'b10001_101010_11100;
end_screen[29][14] = 16'b10001_101010_11100;
end_screen[29][15] = 16'b10001_101010_11100;
end_screen[29][16] = 16'b10001_101010_11100;
end_screen[29][17] = 16'b10001_101010_11100;
end_screen[29][18] = 16'b10001_101010_11100;
end_screen[29][19] = 16'b10001_101010_11100;
end_screen[29][20] = 16'b10001_101010_11100;
end_screen[29][21] = 16'b10001_101010_11100;
end_screen[29][22] = 16'b10001_101010_11100;
end_screen[29][23] = 16'b10001_101010_11100;
end_screen[29][24] = 16'b10010_101000_11001;
end_screen[29][25] = 16'b10011_100010_01111;
end_screen[29][26] = 16'b10101_011100_00110;
end_screen[29][27] = 16'b10011_011000_00100;
end_screen[29][28] = 16'b01111_010010_00010;
end_screen[29][29] = 16'b01100_001100_00001;
end_screen[29][30] = 16'b01010_001010_00000;
end_screen[29][31] = 16'b01010_001000_00000;
end_screen[29][32] = 16'b10000_010100_00100;
end_screen[29][33] = 16'b10110_100000_01001;
end_screen[29][34] = 16'b10010_010111_00100;
end_screen[29][35] = 16'b01111_010111_01000;
end_screen[29][36] = 16'b01111_011000_01001;
end_screen[29][37] = 16'b10000_011010_01010;
end_screen[29][38] = 16'b11111_111111_11111;
end_screen[29][39] = 16'b11111_111111_11111;
end_screen[29][40] = 16'b11111_111111_11111;
end_screen[29][41] = 16'b11111_111111_11111;
end_screen[29][42] = 16'b11111_111111_11111;
end_screen[29][43] = 16'b11111_111111_11111;
end_screen[29][44] = 16'b11111_111111_11111;
end_screen[29][45] = 16'b11111_111111_11111;
end_screen[29][46] = 16'b11111_111111_11111;
end_screen[29][47] = 16'b11111_111111_11111;
end_screen[29][48] = 16'b11111_111111_11111;
end_screen[29][49] = 16'b11111_111111_11111;
end_screen[29][50] = 16'b11111_111111_11111;
end_screen[29][51] = 16'b11111_111111_11111;
end_screen[29][52] = 16'b11111_111111_11111;
end_screen[29][53] = 16'b11111_111111_11111;
end_screen[29][54] = 16'b11111_111111_11111;
end_screen[29][55] = 16'b11111_111111_11111;
end_screen[29][56] = 16'b11111_111111_11111;
end_screen[29][57] = 16'b11111_111111_11111;
end_screen[29][58] = 16'b11111_111111_11111;
end_screen[29][59] = 16'b11000_011011_01000;
end_screen[29][60] = 16'b11001_100000_01010;
end_screen[29][61] = 16'b11001_011111_01001;
end_screen[29][62] = 16'b11011_010111_00011;
end_screen[29][63] = 16'b11011_011000_00100;
end_screen[29][64] = 16'b11011_011000_00011;
end_screen[29][65] = 16'b11011_011000_00100;
end_screen[29][66] = 16'b11011_011000_00100;
end_screen[29][67] = 16'b11011_010111_00011;
end_screen[29][68] = 16'b11010_010010_00010;
end_screen[29][69] = 16'b11010_010100_00010;
end_screen[29][70] = 16'b11011_010101_00010;
end_screen[29][71] = 16'b11100_011110_00110;
end_screen[29][72] = 16'b10111_101010_10100;
end_screen[29][73] = 16'b10011_101011_11011;
end_screen[29][74] = 16'b10001_101010_11100;
end_screen[29][75] = 16'b10001_101010_11100;
end_screen[29][76] = 16'b10001_101010_11100;
end_screen[29][77] = 16'b10001_101010_11100;
end_screen[29][78] = 16'b10001_101010_11100;
end_screen[29][79] = 16'b10001_101010_11100;
end_screen[29][80] = 16'b10001_101010_11100;
end_screen[29][81] = 16'b10001_101010_11100;
end_screen[29][82] = 16'b10001_101010_11100;
end_screen[29][83] = 16'b10001_101010_11100;
end_screen[29][84] = 16'b10001_101010_11100;
end_screen[29][85] = 16'b10001_101010_11100;
end_screen[29][86] = 16'b10001_101010_11100;
end_screen[29][87] = 16'b10001_101010_11100;
end_screen[29][88] = 16'b10001_101010_11100;
end_screen[29][89] = 16'b10001_101010_11100;
end_screen[29][90] = 16'b10001_101010_11100;
end_screen[29][91] = 16'b10001_101010_11100;
end_screen[29][92] = 16'b10001_101010_11100;
end_screen[29][93] = 16'b10001_101010_11100;
end_screen[29][94] = 16'b10001_101010_11100;
end_screen[29][95] = 16'b10001_101010_11100;
end_screen[30][0] = 16'b10001_101010_11100;
end_screen[30][1] = 16'b10001_101010_11100;
end_screen[30][2] = 16'b10001_101010_11100;
end_screen[30][3] = 16'b10001_101010_11100;
end_screen[30][4] = 16'b10001_101010_11100;
end_screen[30][5] = 16'b10001_101010_11100;
end_screen[30][6] = 16'b10001_101010_11100;
end_screen[30][7] = 16'b10001_101010_11100;
end_screen[30][8] = 16'b10001_101010_11100;
end_screen[30][9] = 16'b10001_101010_11100;
end_screen[30][10] = 16'b10001_101010_11100;
end_screen[30][11] = 16'b10001_101010_11100;
end_screen[30][12] = 16'b10001_101010_11100;
end_screen[30][13] = 16'b10001_101010_11100;
end_screen[30][14] = 16'b10001_101010_11100;
end_screen[30][15] = 16'b10001_101010_11100;
end_screen[30][16] = 16'b10001_101010_11100;
end_screen[30][17] = 16'b10001_101010_11100;
end_screen[30][18] = 16'b10001_101010_11100;
end_screen[30][19] = 16'b10001_101010_11100;
end_screen[30][20] = 16'b10001_101010_11100;
end_screen[30][21] = 16'b10001_101010_11100;
end_screen[30][22] = 16'b10001_101010_11100;
end_screen[30][23] = 16'b10001_101010_11100;
end_screen[30][24] = 16'b10010_100011_10010;
end_screen[30][25] = 16'b10010_010110_00011;
end_screen[30][26] = 16'b10111_100000_00111;
end_screen[30][27] = 16'b10000_010011_00011;
end_screen[30][28] = 16'b01010_001010_00000;
end_screen[30][29] = 16'b01011_001010_00000;
end_screen[30][30] = 16'b01100_001100_00001;
end_screen[30][31] = 16'b01101_001101_00000;
end_screen[30][32] = 16'b10100_011100_00110;
end_screen[30][33] = 16'b11011_101011_01101;
end_screen[30][34] = 16'b10101_011101_00110;
end_screen[30][35] = 16'b11111_111111_11111;
end_screen[30][36] = 16'b11111_111111_11111;
end_screen[30][37] = 16'b11111_111111_11111;
end_screen[30][38] = 16'b11111_111111_11111;
end_screen[30][39] = 16'b11111_111111_11111;
end_screen[30][40] = 16'b11111_111111_11111;
end_screen[30][41] = 16'b11111_111111_11111;
end_screen[30][42] = 16'b11111_111111_11111;
end_screen[30][43] = 16'b11111_111111_11111;
end_screen[30][44] = 16'b11111_111111_11111;
end_screen[30][45] = 16'b11111_111111_11111;
end_screen[30][46] = 16'b11111_111111_11111;
end_screen[30][47] = 16'b11111_111111_11111;
end_screen[30][48] = 16'b11111_111111_11111;
end_screen[30][49] = 16'b11111_111111_11111;
end_screen[30][50] = 16'b11111_111111_11111;
end_screen[30][51] = 16'b11111_111111_11111;
end_screen[30][52] = 16'b10100_101001_10100;
end_screen[30][53] = 16'b10100_101001_10100;
end_screen[30][54] = 16'b10100_101001_10100;
end_screen[30][55] = 16'b11111_111111_11111;
end_screen[30][56] = 16'b11111_111111_11111;
end_screen[30][57] = 16'b11111_111111_11111;
end_screen[30][58] = 16'b11111_111111_11111;
end_screen[30][59] = 16'b11111_111111_11111;
end_screen[30][60] = 16'b11111_111111_11111;
end_screen[30][61] = 16'b11111_111111_11111;
end_screen[30][62] = 16'b11011_011000_00100;
end_screen[30][63] = 16'b11100_011001_00100;
end_screen[30][64] = 16'b11011_010111_00011;
end_screen[30][65] = 16'b11100_011001_00100;
end_screen[30][66] = 16'b11100_011001_00100;
end_screen[30][67] = 16'b11011_010111_00011;
end_screen[30][68] = 16'b11010_010011_00010;
end_screen[30][69] = 16'b11010_010101_00010;
end_screen[30][70] = 16'b11011_010110_00011;
end_screen[30][71] = 16'b11011_010001_00001;
end_screen[30][72] = 16'b11011_100100_01010;
end_screen[30][73] = 16'b11011_110010_10001;
end_screen[30][74] = 16'b10111_101101_10100;
end_screen[30][75] = 16'b10001_101010_11100;
end_screen[30][76] = 16'b10001_101010_11100;
end_screen[30][77] = 16'b10001_101010_11100;
end_screen[30][78] = 16'b10001_101010_11100;
end_screen[30][79] = 16'b10001_101010_11100;
end_screen[30][80] = 16'b10001_101010_11100;
end_screen[30][81] = 16'b10001_101010_11100;
end_screen[30][82] = 16'b10001_101010_11100;
end_screen[30][83] = 16'b10001_101010_11100;
end_screen[30][84] = 16'b10001_101010_11100;
end_screen[30][85] = 16'b10001_101010_11100;
end_screen[30][86] = 16'b10001_101010_11100;
end_screen[30][87] = 16'b10001_101010_11100;
end_screen[30][88] = 16'b10001_101010_11100;
end_screen[30][89] = 16'b10001_101010_11100;
end_screen[30][90] = 16'b10001_101010_11100;
end_screen[30][91] = 16'b10001_101010_11100;
end_screen[30][92] = 16'b10001_101010_11100;
end_screen[30][93] = 16'b10001_101010_11100;
end_screen[30][94] = 16'b10001_101010_11100;
end_screen[30][95] = 16'b10001_101010_11100;
end_screen[31][0] = 16'b10001_101010_11100;
end_screen[31][1] = 16'b10001_101010_11100;
end_screen[31][2] = 16'b10001_101010_11100;
end_screen[31][3] = 16'b10001_101010_11100;
end_screen[31][4] = 16'b10001_101010_11100;
end_screen[31][5] = 16'b10001_101010_11100;
end_screen[31][6] = 16'b10001_101010_11100;
end_screen[31][7] = 16'b10001_101010_11100;
end_screen[31][8] = 16'b10001_101010_11100;
end_screen[31][9] = 16'b10001_101010_11100;
end_screen[31][10] = 16'b10001_101010_11100;
end_screen[31][11] = 16'b10001_101010_11100;
end_screen[31][12] = 16'b10001_101010_11100;
end_screen[31][13] = 16'b10001_101010_11100;
end_screen[31][14] = 16'b10001_101010_11100;
end_screen[31][15] = 16'b10001_101010_11100;
end_screen[31][16] = 16'b10001_101010_11100;
end_screen[31][17] = 16'b10001_101010_11100;
end_screen[31][18] = 16'b10001_101010_11100;
end_screen[31][19] = 16'b10001_101010_11100;
end_screen[31][20] = 16'b10001_101010_11100;
end_screen[31][21] = 16'b10001_101010_11100;
end_screen[31][22] = 16'b10001_101010_11100;
end_screen[31][23] = 16'b10001_101010_11100;
end_screen[31][24] = 16'b10010_100011_10011;
end_screen[31][25] = 16'b10010_010101_00011;
end_screen[31][26] = 16'b10011_011001_00100;
end_screen[31][27] = 16'b01011_001100_00001;
end_screen[31][28] = 16'b01011_001011_00001;
end_screen[31][29] = 16'b01011_001011_00001;
end_screen[31][30] = 16'b01101_001101_00001;
end_screen[31][31] = 16'b01111_010001_00010;
end_screen[31][32] = 16'b01111_010001_00010;
end_screen[31][33] = 16'b01110_001111_00001;
end_screen[31][34] = 16'b01100_001100_00001;
end_screen[31][35] = 16'b11111_111111_11111;
end_screen[31][36] = 16'b11111_111111_11111;
end_screen[31][37] = 16'b11111_111111_11111;
end_screen[31][38] = 16'b11111_111111_11111;
end_screen[31][39] = 16'b11111_111111_11111;
end_screen[31][40] = 16'b11111_111111_11111;
end_screen[31][41] = 16'b11111_111111_11111;
end_screen[31][42] = 16'b11111_111111_11111;
end_screen[31][43] = 16'b11111_111111_11111;
end_screen[31][44] = 16'b11111_111111_11111;
end_screen[31][45] = 16'b11111_111111_11111;
end_screen[31][46] = 16'b11111_111111_11111;
end_screen[31][47] = 16'b11111_111111_11111;
end_screen[31][48] = 16'b11111_111111_11111;
end_screen[31][49] = 16'b11111_111111_11111;
end_screen[31][50] = 16'b11111_111111_11111;
end_screen[31][51] = 16'b11111_111111_11111;
end_screen[31][52] = 16'b10100_101001_10100;
end_screen[31][53] = 16'b10100_101001_10100;
end_screen[31][54] = 16'b10100_101001_10100;
end_screen[31][55] = 16'b11111_111111_11111;
end_screen[31][56] = 16'b11111_111111_11111;
end_screen[31][57] = 16'b11111_111111_11111;
end_screen[31][58] = 16'b11111_111111_11111;
end_screen[31][59] = 16'b11111_111111_11111;
end_screen[31][60] = 16'b11111_111111_11111;
end_screen[31][61] = 16'b11111_111111_11111;
end_screen[31][62] = 16'b11011_010101_00011;
end_screen[31][63] = 16'b11011_010101_00011;
end_screen[31][64] = 16'b11011_011000_00100;
end_screen[31][65] = 16'b11011_011000_00100;
end_screen[31][66] = 16'b11011_010110_00011;
end_screen[31][67] = 16'b11011_010111_00011;
end_screen[31][68] = 16'b11011_011000_00100;
end_screen[31][69] = 16'b11011_011000_00100;
end_screen[31][70] = 16'b11010_010010_00010;
end_screen[31][71] = 16'b11010_001111_00000;
end_screen[31][72] = 16'b11011_100011_01010;
end_screen[31][73] = 16'b11011_110001_10000;
end_screen[31][74] = 16'b11100_110000_10000;
end_screen[31][75] = 16'b10111_101110_10101;
end_screen[31][76] = 16'b10001_101010_11100;
end_screen[31][77] = 16'b10001_101010_11100;
end_screen[31][78] = 16'b10001_101010_11100;
end_screen[31][79] = 16'b10001_101010_11100;
end_screen[31][80] = 16'b10001_101010_11100;
end_screen[31][81] = 16'b10001_101010_11100;
end_screen[31][82] = 16'b10001_101010_11100;
end_screen[31][83] = 16'b10001_101010_11100;
end_screen[31][84] = 16'b10001_101010_11100;
end_screen[31][85] = 16'b10001_101010_11100;
end_screen[31][86] = 16'b10001_101010_11100;
end_screen[31][87] = 16'b10001_101010_11100;
end_screen[31][88] = 16'b10001_101010_11100;
end_screen[31][89] = 16'b10001_101010_11100;
end_screen[31][90] = 16'b10001_101010_11100;
end_screen[31][91] = 16'b10001_101010_11100;
end_screen[31][92] = 16'b10001_101010_11100;
end_screen[31][93] = 16'b10001_101010_11100;
end_screen[31][94] = 16'b10001_101010_11100;
end_screen[31][95] = 16'b10001_101010_11100;
end_screen[32][0] = 16'b10001_101010_11100;
end_screen[32][1] = 16'b10001_101010_11100;
end_screen[32][2] = 16'b10001_101010_11100;
end_screen[32][3] = 16'b10001_101010_11100;
end_screen[32][4] = 16'b10001_101010_11100;
end_screen[32][5] = 16'b10001_101010_11100;
end_screen[32][6] = 16'b10001_101010_11100;
end_screen[32][7] = 16'b10001_101010_11100;
end_screen[32][8] = 16'b10001_101010_11100;
end_screen[32][9] = 16'b10001_101010_11100;
end_screen[32][10] = 16'b10001_101010_11100;
end_screen[32][11] = 16'b10001_101010_11100;
end_screen[32][12] = 16'b10001_101010_11100;
end_screen[32][13] = 16'b10001_101010_11100;
end_screen[32][14] = 16'b10001_101010_11100;
end_screen[32][15] = 16'b10001_101010_11100;
end_screen[32][16] = 16'b10001_101010_11100;
end_screen[32][17] = 16'b10001_101010_11100;
end_screen[32][18] = 16'b10001_101010_11100;
end_screen[32][19] = 16'b10001_101010_11100;
end_screen[32][20] = 16'b10001_101010_11100;
end_screen[32][21] = 16'b10001_101010_11100;
end_screen[32][22] = 16'b01101_100000_10000;
end_screen[32][23] = 16'b01110_011111_01110;
end_screen[32][24] = 16'b01101_011011_01010;
end_screen[32][25] = 16'b01101_010101_00011;
end_screen[32][26] = 16'b01111_010110_00100;
end_screen[32][27] = 16'b01011_001011_00001;
end_screen[32][28] = 16'b01011_001011_00001;
end_screen[32][29] = 16'b01100_001100_00001;
end_screen[32][30] = 16'b01110_010000_00010;
end_screen[32][31] = 16'b01111_010001_00010;
end_screen[32][32] = 16'b01101_001110_00001;
end_screen[32][33] = 16'b01011_001011_00000;
end_screen[32][34] = 16'b01100_001100_00001;
end_screen[32][35] = 16'b11111_111111_11111;
end_screen[32][36] = 16'b11111_111111_11111;
end_screen[32][37] = 16'b11111_111111_11111;
end_screen[32][38] = 16'b11111_111111_11111;
end_screen[32][39] = 16'b11111_111111_11111;
end_screen[32][40] = 16'b11111_111111_11111;
end_screen[32][41] = 16'b11111_111111_11111;
end_screen[32][42] = 16'b11111_111111_11111;
end_screen[32][43] = 16'b11111_111111_11111;
end_screen[32][44] = 16'b11111_111111_11111;
end_screen[32][45] = 16'b11111_111111_11111;
end_screen[32][46] = 16'b11111_111111_11111;
end_screen[32][47] = 16'b11111_111111_11111;
end_screen[32][48] = 16'b11111_111111_11111;
end_screen[32][49] = 16'b11111_111111_11111;
end_screen[32][50] = 16'b11111_111111_11111;
end_screen[32][51] = 16'b11111_111111_11111;
end_screen[32][52] = 16'b10100_101001_10100;
end_screen[32][53] = 16'b10100_101001_10100;
end_screen[32][54] = 16'b10100_101001_10100;
end_screen[32][55] = 16'b11111_111111_11111;
end_screen[32][56] = 16'b11111_111111_11111;
end_screen[32][57] = 16'b11111_111111_11111;
end_screen[32][58] = 16'b11111_111111_11111;
end_screen[32][59] = 16'b11111_111111_11111;
end_screen[32][60] = 16'b11111_111111_11111;
end_screen[32][61] = 16'b11111_111111_11111;
end_screen[32][62] = 16'b11011_010101_00011;
end_screen[32][63] = 16'b11011_010111_00011;
end_screen[32][64] = 16'b11011_011001_00100;
end_screen[32][65] = 16'b11011_010101_00011;
end_screen[32][66] = 16'b11011_010111_00011;
end_screen[32][67] = 16'b11010_010101_00010;
end_screen[32][68] = 16'b11010_010100_00010;
end_screen[32][69] = 16'b11011_010110_00011;
end_screen[32][70] = 16'b11011_010110_00011;
end_screen[32][71] = 16'b11010_010011_00010;
end_screen[32][72] = 16'b11011_011010_00101;
end_screen[32][73] = 16'b11100_101011_01101;
end_screen[32][74] = 16'b11100_110010_10010;
end_screen[32][75] = 16'b11011_101110_01111;
end_screen[32][76] = 16'b11000_101101_10100;
end_screen[32][77] = 16'b10001_101010_11100;
end_screen[32][78] = 16'b10001_101010_11100;
end_screen[32][79] = 16'b10001_101010_11100;
end_screen[32][80] = 16'b10001_101010_11100;
end_screen[32][81] = 16'b10001_101010_11100;
end_screen[32][82] = 16'b10001_101010_11100;
end_screen[32][83] = 16'b10001_101010_11100;
end_screen[32][84] = 16'b10001_101010_11100;
end_screen[32][85] = 16'b10001_101010_11100;
end_screen[32][86] = 16'b10001_101010_11100;
end_screen[32][87] = 16'b10001_101010_11100;
end_screen[32][88] = 16'b10001_101010_11100;
end_screen[32][89] = 16'b10001_101010_11100;
end_screen[32][90] = 16'b10001_101010_11100;
end_screen[32][91] = 16'b10001_101010_11100;
end_screen[32][92] = 16'b10001_101010_11100;
end_screen[32][93] = 16'b10001_101010_11100;
end_screen[32][94] = 16'b10001_101010_11100;
end_screen[32][95] = 16'b10001_101010_11100;
end_screen[33][0] = 16'b10001_101010_11100;
end_screen[33][1] = 16'b10001_101010_11100;
end_screen[33][2] = 16'b10001_101010_11100;
end_screen[33][3] = 16'b10001_101010_11100;
end_screen[33][4] = 16'b10001_101010_11100;
end_screen[33][5] = 16'b10001_101010_11100;
end_screen[33][6] = 16'b10001_101010_11100;
end_screen[33][7] = 16'b10001_101010_11100;
end_screen[33][8] = 16'b10001_101010_11100;
end_screen[33][9] = 16'b10001_101010_11100;
end_screen[33][10] = 16'b10001_101010_11100;
end_screen[33][11] = 16'b10001_101010_11100;
end_screen[33][12] = 16'b10001_101010_11100;
end_screen[33][13] = 16'b10001_101010_11100;
end_screen[33][14] = 16'b10001_101010_11100;
end_screen[33][15] = 16'b10001_101010_11100;
end_screen[33][16] = 16'b10001_101010_11100;
end_screen[33][17] = 16'b10001_101010_11100;
end_screen[33][18] = 16'b10001_101010_11100;
end_screen[33][19] = 16'b10001_101010_11100;
end_screen[33][20] = 16'b10001_101010_11100;
end_screen[33][21] = 16'b01111_100011_10011;
end_screen[33][22] = 16'b01101_011011_00101;
end_screen[33][23] = 16'b01111_011110_00111;
end_screen[33][24] = 16'b10010_100011_01001;
end_screen[33][25] = 16'b10000_011111_01000;
end_screen[33][26] = 16'b01100_011001_00101;
end_screen[33][27] = 16'b01100_010011_00011;
end_screen[33][28] = 16'b01100_010010_00011;
end_screen[33][29] = 16'b01100_001100_00000;
end_screen[33][30] = 16'b10101_011101_00111;
end_screen[33][31] = 16'b11001_100100_01000;
end_screen[33][32] = 16'b10001_010101_00011;
end_screen[33][33] = 16'b01010_001001_00000;
end_screen[33][34] = 16'b01100_001100_00001;
end_screen[33][35] = 16'b11111_111111_11111;
end_screen[33][36] = 16'b11111_111111_11111;
end_screen[33][37] = 16'b11111_111111_11111;
end_screen[33][38] = 16'b11111_111111_11111;
end_screen[33][39] = 16'b10100_101001_10100;
end_screen[33][40] = 16'b10100_101001_10100;
end_screen[33][41] = 16'b11111_111111_11111;
end_screen[33][42] = 16'b11111_111111_11111;
end_screen[33][43] = 16'b11111_111111_11111;
end_screen[33][44] = 16'b11111_111111_11111;
end_screen[33][45] = 16'b10100_101001_10100;
end_screen[33][46] = 16'b10100_101001_10100;
end_screen[33][47] = 16'b10100_101001_10100;
end_screen[33][48] = 16'b11111_111111_11111;
end_screen[33][49] = 16'b11111_111111_11111;
end_screen[33][50] = 16'b11111_111111_11111;
end_screen[33][51] = 16'b11111_111111_11111;
end_screen[33][52] = 16'b10100_101001_10100;
end_screen[33][53] = 16'b10100_101001_10100;
end_screen[33][54] = 16'b10100_101001_10100;
end_screen[33][55] = 16'b11111_111111_11111;
end_screen[33][56] = 16'b11111_111111_11111;
end_screen[33][57] = 16'b11111_111111_11111;
end_screen[33][58] = 16'b11111_111111_11111;
end_screen[33][59] = 16'b11111_111111_11111;
end_screen[33][60] = 16'b11111_111111_11111;
end_screen[33][61] = 16'b11111_111111_11111;
end_screen[33][62] = 16'b11011_010110_00011;
end_screen[33][63] = 16'b11100_011011_00101;
end_screen[33][64] = 16'b11100_011001_00100;
end_screen[33][65] = 16'b11011_011000_00100;
end_screen[33][66] = 16'b11011_010111_00011;
end_screen[33][67] = 16'b11010_010010_00010;
end_screen[33][68] = 16'b11010_010011_00010;
end_screen[33][69] = 16'b11011_010110_00011;
end_screen[33][70] = 16'b11011_011000_00100;
end_screen[33][71] = 16'b11010_010100_00010;
end_screen[33][72] = 16'b11010_011000_00101;
end_screen[33][73] = 16'b11100_110000_10010;
end_screen[33][74] = 16'b11100_110011_10011;
end_screen[33][75] = 16'b11011_110001_10010;
end_screen[33][76] = 16'b11100_110010_10011;
end_screen[33][77] = 16'b11011_110001_10011;
end_screen[33][78] = 16'b11010_110000_10100;
end_screen[33][79] = 16'b11010_110001_10100;
end_screen[33][80] = 16'b11010_110000_10100;
end_screen[33][81] = 16'b11010_110001_10100;
end_screen[33][82] = 16'b11010_110000_10100;
end_screen[33][83] = 16'b11010_101111_10011;
end_screen[33][84] = 16'b11010_110000_10100;
end_screen[33][85] = 16'b11010_110000_10100;
end_screen[33][86] = 16'b10101_101101_11001;
end_screen[33][87] = 16'b10001_101010_11100;
end_screen[33][88] = 16'b10001_101010_11100;
end_screen[33][89] = 16'b10001_101010_11100;
end_screen[33][90] = 16'b10001_101010_11100;
end_screen[33][91] = 16'b10001_101010_11100;
end_screen[33][92] = 16'b10001_101010_11100;
end_screen[33][93] = 16'b10001_101010_11100;
end_screen[33][94] = 16'b10001_101010_11100;
end_screen[33][95] = 16'b10001_101010_11100;
end_screen[34][0] = 16'b10001_101010_11100;
end_screen[34][1] = 16'b10001_101010_11100;
end_screen[34][2] = 16'b10001_101010_11100;
end_screen[34][3] = 16'b10001_101010_11100;
end_screen[34][4] = 16'b10001_101010_11100;
end_screen[34][5] = 16'b10001_101010_11100;
end_screen[34][6] = 16'b10001_101010_11100;
end_screen[34][7] = 16'b10001_101010_11100;
end_screen[34][8] = 16'b10001_101010_11100;
end_screen[34][9] = 16'b10001_101010_11100;
end_screen[34][10] = 16'b10001_101010_11100;
end_screen[34][11] = 16'b10001_101010_11100;
end_screen[34][12] = 16'b10011_101100_11010;
end_screen[34][13] = 16'b10011_101100_11010;
end_screen[34][14] = 16'b10011_101100_11010;
end_screen[34][15] = 16'b10011_101100_11010;
end_screen[34][16] = 16'b10011_101011_11010;
end_screen[34][17] = 16'b10011_101011_11010;
end_screen[34][18] = 16'b10011_101100_11010;
end_screen[34][19] = 16'b10011_101011_11001;
end_screen[34][20] = 16'b10000_100110_10110;
end_screen[34][21] = 16'b01100_011001_00101;
end_screen[34][22] = 16'b01111_011111_00111;
end_screen[34][23] = 16'b10010_100101_01010;
end_screen[34][24] = 16'b10111_101100_01110;
end_screen[34][25] = 16'b10010_100011_01010;
end_screen[34][26] = 16'b01100_011011_00101;
end_screen[34][27] = 16'b10000_100000_00111;
end_screen[34][28] = 16'b01110_011110_00111;
end_screen[34][29] = 16'b01100_010001_00010;
end_screen[34][30] = 16'b01111_010001_00010;
end_screen[34][31] = 16'b10000_010011_00011;
end_screen[34][32] = 16'b01101_001110_00001;
end_screen[34][33] = 16'b01011_001011_00001;
end_screen[34][34] = 16'b01100_001100_00001;
end_screen[34][35] = 16'b11111_111111_11111;
end_screen[34][36] = 16'b11111_111111_11111;
end_screen[34][37] = 16'b11111_111111_11111;
end_screen[34][38] = 16'b11111_111111_11111;
end_screen[34][39] = 16'b10100_101001_10100;
end_screen[34][40] = 16'b10100_101001_10100;
end_screen[34][41] = 16'b11111_111111_11111;
end_screen[34][42] = 16'b11111_111111_11111;
end_screen[34][43] = 16'b11111_111111_11111;
end_screen[34][44] = 16'b11111_111111_11111;
end_screen[34][45] = 16'b10100_101001_10100;
end_screen[34][46] = 16'b10100_101001_10100;
end_screen[34][47] = 16'b10100_101001_10100;
end_screen[34][48] = 16'b11111_111111_11111;
end_screen[34][49] = 16'b11111_111111_11111;
end_screen[34][50] = 16'b11111_111111_11111;
end_screen[34][51] = 16'b11111_111111_11111;
end_screen[34][52] = 16'b10100_101001_10100;
end_screen[34][53] = 16'b10100_101001_10100;
end_screen[34][54] = 16'b10100_101001_10100;
end_screen[34][55] = 16'b11111_111111_11111;
end_screen[34][56] = 16'b11111_111111_11111;
end_screen[34][57] = 16'b11111_111111_11111;
end_screen[34][58] = 16'b11111_111111_11111;
end_screen[34][59] = 16'b11111_111111_11111;
end_screen[34][60] = 16'b11111_111111_11111;
end_screen[34][61] = 16'b11111_111111_11111;
end_screen[34][62] = 16'b11011_010101_00011;
end_screen[34][63] = 16'b11011_010111_00011;
end_screen[34][64] = 16'b11010_010101_00011;
end_screen[34][65] = 16'b11010_010011_00010;
end_screen[34][66] = 16'b11010_010100_00010;
end_screen[34][67] = 16'b11010_010100_00010;
end_screen[34][68] = 16'b11011_010110_00011;
end_screen[34][69] = 16'b11011_100100_01011;
end_screen[34][70] = 16'b11011_101011_01111;
end_screen[34][71] = 16'b11011_101011_10000;
end_screen[34][72] = 16'b11100_101110_10001;
end_screen[34][73] = 16'b11011_110000_10010;
end_screen[34][74] = 16'b11010_101011_01110;
end_screen[34][75] = 16'b11001_101011_01110;
end_screen[34][76] = 16'b11001_101011_01110;
end_screen[34][77] = 16'b11001_101011_01110;
end_screen[34][78] = 16'b11001_101011_01110;
end_screen[34][79] = 16'b11001_101011_01110;
end_screen[34][80] = 16'b11001_101011_01110;
end_screen[34][81] = 16'b11001_101011_01110;
end_screen[34][82] = 16'b11001_101010_01110;
end_screen[34][83] = 16'b11001_101010_01110;
end_screen[34][84] = 16'b11001_101010_01110;
end_screen[34][85] = 16'b11010_101101_10000;
end_screen[34][86] = 16'b11011_110000_10011;
end_screen[34][87] = 16'b11001_110000_10101;
end_screen[34][88] = 16'b11001_110000_10101;
end_screen[34][89] = 16'b10111_101110_10110;
end_screen[34][90] = 16'b10001_101010_11100;
end_screen[34][91] = 16'b10001_101010_11100;
end_screen[34][92] = 16'b10001_101010_11100;
end_screen[34][93] = 16'b10001_101010_11100;
end_screen[34][94] = 16'b10001_101010_11100;
end_screen[34][95] = 16'b10001_101010_11100;
end_screen[35][0] = 16'b10001_101010_11100;
end_screen[35][1] = 16'b10001_101010_11100;
end_screen[35][2] = 16'b10001_101010_11100;
end_screen[35][3] = 16'b10001_101010_11100;
end_screen[35][4] = 16'b10001_101010_11100;
end_screen[35][5] = 16'b10001_101010_11100;
end_screen[35][6] = 16'b10001_101010_11100;
end_screen[35][7] = 16'b10001_101010_11100;
end_screen[35][8] = 16'b10010_101010_11011;
end_screen[35][9] = 16'b10010_101011_11011;
end_screen[35][10] = 16'b10010_101011_11011;
end_screen[35][11] = 16'b10101_101100_10111;
end_screen[35][12] = 16'b11011_101111_10000;
end_screen[35][13] = 16'b11100_110001_10001;
end_screen[35][14] = 16'b11100_110001_10001;
end_screen[35][15] = 16'b11011_110000_10000;
end_screen[35][16] = 16'b11011_101111_01111;
end_screen[35][17] = 16'b11011_101110_01111;
end_screen[35][18] = 16'b11100_101111_10000;
end_screen[35][19] = 16'b10111_101001_01100;
end_screen[35][20] = 16'b01110_011101_00110;
end_screen[35][21] = 16'b01111_100000_00111;
end_screen[35][22] = 16'b01111_011111_00111;
end_screen[35][23] = 16'b10001_100011_01001;
end_screen[35][24] = 16'b10001_100011_01001;
end_screen[35][25] = 16'b10000_100001_01000;
end_screen[35][26] = 16'b10001_100010_01001;
end_screen[35][27] = 16'b10010_100101_01010;
end_screen[35][28] = 16'b10010_100100_01010;
end_screen[35][29] = 16'b01101_011011_00110;
end_screen[35][30] = 16'b01011_001110_00010;
end_screen[35][31] = 16'b01010_001010_00000;
end_screen[35][32] = 16'b01010_001001_00000;
end_screen[35][33] = 16'b01011_001100_00001;
end_screen[35][34] = 16'b01110_001111_00001;
end_screen[35][35] = 16'b11111_111111_11111;
end_screen[35][36] = 16'b11111_111111_11111;
end_screen[35][37] = 16'b11111_111111_11111;
end_screen[35][38] = 16'b11111_111111_11111;
end_screen[35][39] = 16'b10100_101001_10100;
end_screen[35][40] = 16'b10100_101001_10100;
end_screen[35][41] = 16'b11111_111111_11111;
end_screen[35][42] = 16'b11111_111111_11111;
end_screen[35][43] = 16'b11111_111111_11111;
end_screen[35][44] = 16'b11111_111111_11111;
end_screen[35][45] = 16'b10100_101001_10100;
end_screen[35][46] = 16'b10100_101001_10100;
end_screen[35][47] = 16'b10100_101001_10100;
end_screen[35][48] = 16'b11111_111111_11111;
end_screen[35][49] = 16'b11111_111111_11111;
end_screen[35][50] = 16'b11111_111111_11111;
end_screen[35][51] = 16'b11111_111111_11111;
end_screen[35][52] = 16'b10100_101001_10100;
end_screen[35][53] = 16'b10100_101001_10100;
end_screen[35][54] = 16'b10100_101001_10100;
end_screen[35][55] = 16'b11111_111111_11111;
end_screen[35][56] = 16'b11111_111111_11111;
end_screen[35][57] = 16'b11111_111111_11111;
end_screen[35][58] = 16'b11111_111111_11111;
end_screen[35][59] = 16'b11111_111111_11111;
end_screen[35][60] = 16'b11111_111111_11111;
end_screen[35][61] = 16'b11111_111111_11111;
end_screen[35][62] = 16'b11010_010100_00010;
end_screen[35][63] = 16'b11011_010110_00011;
end_screen[35][64] = 16'b11010_010100_00010;
end_screen[35][65] = 16'b11010_010011_00010;
end_screen[35][66] = 16'b11010_010010_00010;
end_screen[35][67] = 16'b11010_010101_00010;
end_screen[35][68] = 16'b11011_100101_01100;
end_screen[35][69] = 16'b11011_110000_10010;
end_screen[35][70] = 16'b11010_101110_10000;
end_screen[35][71] = 16'b11010_101011_01110;
end_screen[35][72] = 16'b11010_101010_01110;
end_screen[35][73] = 16'b11001_101011_01110;
end_screen[35][74] = 16'b11001_101011_01101;
end_screen[35][75] = 16'b11001_101100_01110;
end_screen[35][76] = 16'b11001_101100_01101;
end_screen[35][77] = 16'b11001_101100_01110;
end_screen[35][78] = 16'b11001_101100_01110;
end_screen[35][79] = 16'b11001_101100_01101;
end_screen[35][80] = 16'b11001_101100_01101;
end_screen[35][81] = 16'b11001_101100_01101;
end_screen[35][82] = 16'b11001_101100_01110;
end_screen[35][83] = 16'b11001_101100_01110;
end_screen[35][84] = 16'b11001_101011_01101;
end_screen[35][85] = 16'b11001_101010_01101;
end_screen[35][86] = 16'b11001_101010_01110;
end_screen[35][87] = 16'b11010_101101_10000;
end_screen[35][88] = 16'b11011_101111_10001;
end_screen[35][89] = 16'b11011_110000_10010;
end_screen[35][90] = 16'b11000_101110_10101;
end_screen[35][91] = 16'b10001_101010_11100;
end_screen[35][92] = 16'b10001_101010_11100;
end_screen[35][93] = 16'b10001_101010_11100;
end_screen[35][94] = 16'b10001_101010_11100;
end_screen[35][95] = 16'b10001_101010_11100;
end_screen[36][0] = 16'b10001_101010_11100;
end_screen[36][1] = 16'b10001_101010_11100;
end_screen[36][2] = 16'b10001_101010_11100;
end_screen[36][3] = 16'b10001_101010_11100;
end_screen[36][4] = 16'b10001_101010_11100;
end_screen[36][5] = 16'b10001_101010_11100;
end_screen[36][6] = 16'b10001_101010_11100;
end_screen[36][7] = 16'b10001_101010_11100;
end_screen[36][8] = 16'b11000_101101_10011;
end_screen[36][9] = 16'b11100_110000_10000;
end_screen[36][10] = 16'b11011_101111_10000;
end_screen[36][11] = 16'b11011_101110_01111;
end_screen[36][12] = 16'b11011_101110_01111;
end_screen[36][13] = 16'b11011_101101_01110;
end_screen[36][14] = 16'b11011_101100_01110;
end_screen[36][15] = 16'b11011_101100_01110;
end_screen[36][16] = 16'b11010_101011_01110;
end_screen[36][17] = 16'b11100_101110_01111;
end_screen[36][18] = 16'b10111_101001_01100;
end_screen[36][19] = 16'b01111_100000_00111;
end_screen[36][20] = 16'b10010_100100_01001;
end_screen[36][21] = 16'b10010_100100_01001;
end_screen[36][22] = 16'b10000_100001_01000;
end_screen[36][23] = 16'b01111_011111_00111;
end_screen[36][24] = 16'b10010_100100_01010;
end_screen[36][25] = 16'b10011_100110_01010;
end_screen[36][26] = 16'b10001_100011_01001;
end_screen[36][27] = 16'b10011_100110_01011;
end_screen[36][28] = 16'b10000_100000_01000;
end_screen[36][29] = 16'b01101_011100_00110;
end_screen[36][30] = 16'b01101_011011_00101;
end_screen[36][31] = 16'b01101_010100_00011;
end_screen[36][32] = 16'b01110_001111_00001;
end_screen[36][33] = 16'b01100_001100_00001;
end_screen[36][34] = 16'b01011_001011_00001;
end_screen[36][35] = 16'b01011_001100_00001;
end_screen[36][36] = 16'b01010_001010_00001;
end_screen[36][37] = 16'b01001_001001_00000;
end_screen[36][38] = 16'b01001_001001_00000;
end_screen[36][39] = 16'b10100_101001_10100;
end_screen[36][40] = 16'b10100_101001_10100;
end_screen[36][41] = 16'b11111_111111_11111;
end_screen[36][42] = 16'b11111_111111_11111;
end_screen[36][43] = 16'b11111_111111_11111;
end_screen[36][44] = 16'b11111_111111_11111;
end_screen[36][45] = 16'b10100_101001_10100;
end_screen[36][46] = 16'b10100_101001_10100;
end_screen[36][47] = 16'b10100_101001_10100;
end_screen[36][48] = 16'b11111_111111_11111;
end_screen[36][49] = 16'b11111_111111_11111;
end_screen[36][50] = 16'b11111_111111_11111;
end_screen[36][51] = 16'b11111_111111_11111;
end_screen[36][52] = 16'b10100_101001_10100;
end_screen[36][53] = 16'b10100_101001_10100;
end_screen[36][54] = 16'b10100_101001_10100;
end_screen[36][55] = 16'b11111_111111_11111;
end_screen[36][56] = 16'b11111_111111_11111;
end_screen[36][57] = 16'b11111_111111_11111;
end_screen[36][58] = 16'b11001_010100_00011;
end_screen[36][59] = 16'b11001_010100_00011;
end_screen[36][60] = 16'b11001_010011_00011;
end_screen[36][61] = 16'b11001_010011_00011;
end_screen[36][62] = 16'b11010_010101_00010;
end_screen[36][63] = 16'b11010_010011_00010;
end_screen[36][64] = 16'b11011_010101_00011;
end_screen[36][65] = 16'b11011_010110_00011;
end_screen[36][66] = 16'b11010_010100_00010;
end_screen[36][67] = 16'b11011_100101_01100;
end_screen[36][68] = 16'b11010_101100_01111;
end_screen[36][69] = 16'b11001_101010_01101;
end_screen[36][70] = 16'b11001_101011_01110;
end_screen[36][71] = 16'b11001_101100_01110;
end_screen[36][72] = 16'b11001_101111_01111;
end_screen[36][73] = 16'b11001_101010_01101;
end_screen[36][74] = 16'b11000_011100_00111;
end_screen[36][75] = 16'b11000_011000_00110;
end_screen[36][76] = 16'b11000_011000_00110;
end_screen[36][77] = 16'b11000_011000_00110;
end_screen[36][78] = 16'b11000_011000_00110;
end_screen[36][79] = 16'b11000_010111_00110;
end_screen[36][80] = 16'b11000_011000_00110;
end_screen[36][81] = 16'b11001_011001_00110;
end_screen[36][82] = 16'b11001_011001_00110;
end_screen[36][83] = 16'b11000_011001_00110;
end_screen[36][84] = 16'b11000_011100_00111;
end_screen[36][85] = 16'b11001_101001_01100;
end_screen[36][86] = 16'b11001_110000_01111;
end_screen[36][87] = 16'b11001_101110_01111;
end_screen[36][88] = 16'b11010_101101_01111;
end_screen[36][89] = 16'b11010_101011_01110;
end_screen[36][90] = 16'b11010_101011_01110;
end_screen[36][91] = 16'b11000_101111_10110;
end_screen[36][92] = 16'b10001_101010_11100;
end_screen[36][93] = 16'b10001_101010_11100;
end_screen[36][94] = 16'b10001_101010_11100;
end_screen[36][95] = 16'b10001_101010_11100;
end_screen[37][0] = 16'b10001_101010_11100;
end_screen[37][1] = 16'b10001_101010_11100;
end_screen[37][2] = 16'b10001_101010_11100;
end_screen[37][3] = 16'b10001_101010_11100;
end_screen[37][4] = 16'b10001_101010_11100;
end_screen[37][5] = 16'b10001_101010_11100;
end_screen[37][6] = 16'b10001_101010_11100;
end_screen[37][7] = 16'b11000_101100_10010;
end_screen[37][8] = 16'b11011_101100_01110;
end_screen[37][9] = 16'b11011_101111_10000;
end_screen[37][10] = 16'b11011_101010_01011;
end_screen[37][11] = 16'b11011_100100_00101;
end_screen[37][12] = 16'b11011_100100_00101;
end_screen[37][13] = 16'b11010_100001_00011;
end_screen[37][14] = 16'b11001_011110_00010;
end_screen[37][15] = 16'b11001_011111_00011;
end_screen[37][16] = 16'b11001_100100_01000;
end_screen[37][17] = 16'b11100_101101_01111;
end_screen[37][18] = 16'b10110_100110_01011;
end_screen[37][19] = 16'b10000_100001_01000;
end_screen[37][20] = 16'b11100_110100_10011;
end_screen[37][21] = 16'b11101_110110_10100;
end_screen[37][22] = 16'b11100_110011_10011;
end_screen[37][23] = 16'b11010_110001_10001;
end_screen[37][24] = 16'b11100_110011_10011;
end_screen[37][25] = 16'b10110_101011_01110;
end_screen[37][26] = 16'b10000_100001_01000;
end_screen[37][27] = 16'b10001_100011_01001;
end_screen[37][28] = 16'b10000_100001_01000;
end_screen[37][29] = 16'b10011_100101_01010;
end_screen[37][30] = 16'b01101_011100_00110;
end_screen[37][31] = 16'b01111_010110_00100;
end_screen[37][32] = 16'b10000_010010_00010;
end_screen[37][33] = 16'b01111_010001_00010;
end_screen[37][34] = 16'b01110_001111_00010;
end_screen[37][35] = 16'b01101_001110_00001;
end_screen[37][36] = 16'b01101_001110_00001;
end_screen[37][37] = 16'b01101_001111_00001;
end_screen[37][38] = 16'b01101_001111_00001;
end_screen[37][39] = 16'b10100_101001_10100;
end_screen[37][40] = 16'b10100_101001_10100;
end_screen[37][41] = 16'b11111_111111_11111;
end_screen[37][42] = 16'b11111_111111_11111;
end_screen[37][43] = 16'b11111_111111_11111;
end_screen[37][44] = 16'b11111_111111_11111;
end_screen[37][45] = 16'b10100_101001_10100;
end_screen[37][46] = 16'b10100_101001_10100;
end_screen[37][47] = 16'b10100_101001_10100;
end_screen[37][48] = 16'b11111_111111_11111;
end_screen[37][49] = 16'b11111_111111_11111;
end_screen[37][50] = 16'b11111_111111_11111;
end_screen[37][51] = 16'b11111_111111_11111;
end_screen[37][52] = 16'b10100_101001_10100;
end_screen[37][53] = 16'b10100_101001_10100;
end_screen[37][54] = 16'b10100_101001_10100;
end_screen[37][55] = 16'b11111_111111_11111;
end_screen[37][56] = 16'b11111_111111_11111;
end_screen[37][57] = 16'b11111_111111_11111;
end_screen[37][58] = 16'b11010_010011_00010;
end_screen[37][59] = 16'b11010_010011_00010;
end_screen[37][60] = 16'b11010_010011_00010;
end_screen[37][61] = 16'b11011_010110_00011;
end_screen[37][62] = 16'b11011_010110_00011;
end_screen[37][63] = 16'b11010_010011_00010;
end_screen[37][64] = 16'b11001_010010_00010;
end_screen[37][65] = 16'b11010_010100_00011;
end_screen[37][66] = 16'b11011_100100_01011;
end_screen[37][67] = 16'b11010_101100_01111;
end_screen[37][68] = 16'b11001_101010_01110;
end_screen[37][69] = 16'b11001_101110_01110;
end_screen[37][70] = 16'b11001_100110_01011;
end_screen[37][71] = 16'b11000_011100_00111;
end_screen[37][72] = 16'b11000_011101_01000;
end_screen[37][73] = 16'b11000_011000_00110;
end_screen[37][74] = 16'b10110_001001_00000;
end_screen[37][75] = 16'b10110_000110_00000;
end_screen[37][76] = 16'b10111_000110_00000;
end_screen[37][77] = 16'b10111_000110_00000;
end_screen[37][78] = 16'b10111_000111_00000;
end_screen[37][79] = 16'b11000_001000_00000;
end_screen[37][80] = 16'b11000_001001_00000;
end_screen[37][81] = 16'b11000_001001_00000;
end_screen[37][82] = 16'b11000_001001_00000;
end_screen[37][83] = 16'b11001_000110_00000;
end_screen[37][84] = 16'b11001_001000_00000;
end_screen[37][85] = 16'b11001_010110_00101;
end_screen[37][86] = 16'b11000_011110_01000;
end_screen[37][87] = 16'b11000_011100_00111;
end_screen[37][88] = 16'b11001_100100_01010;
end_screen[37][89] = 16'b11001_101101_01110;
end_screen[37][90] = 16'b11001_101011_01110;
end_screen[37][91] = 16'b11001_101010_01110;
end_screen[37][92] = 16'b11000_101111_10110;
end_screen[37][93] = 16'b10010_101011_11011;
end_screen[37][94] = 16'b10001_101010_11100;
end_screen[37][95] = 16'b10001_101010_11100;
end_screen[38][0] = 16'b10001_101010_11100;
end_screen[38][1] = 16'b10001_101010_11100;
end_screen[38][2] = 16'b10001_101010_11100;
end_screen[38][3] = 16'b10001_101010_11100;
end_screen[38][4] = 16'b10010_101011_11011;
end_screen[38][5] = 16'b11010_110000_10011;
end_screen[38][6] = 16'b11010_110000_10100;
end_screen[38][7] = 16'b11100_101111_01111;
end_screen[38][8] = 16'b11011_101110_01111;
end_screen[38][9] = 16'b11010_100110_01001;
end_screen[38][10] = 16'b11011_100011_00100;
end_screen[38][11] = 16'b11100_101000_00111;
end_screen[38][12] = 16'b11101_101011_01001;
end_screen[38][13] = 16'b11100_101010_01001;
end_screen[38][14] = 16'b11010_100100_00110;
end_screen[38][15] = 16'b11001_100101_01000;
end_screen[38][16] = 16'b11001_100001_00101;
end_screen[38][17] = 16'b11000_100000_00101;
end_screen[38][18] = 16'b11001_101010_01101;
end_screen[38][19] = 16'b11011_110100_10011;
end_screen[38][20] = 16'b11111_111000_10110;
end_screen[38][21] = 16'b11111_111001_10111;
end_screen[38][22] = 16'b11111_111001_10110;
end_screen[38][23] = 16'b11110_110111_10101;
end_screen[38][24] = 16'b11110_110111_10101;
end_screen[38][25] = 16'b11101_110101_10100;
end_screen[38][26] = 16'b11011_110001_10010;
end_screen[38][27] = 16'b11000_101101_01111;
end_screen[38][28] = 16'b10011_100101_01010;
end_screen[38][29] = 16'b10001_100010_01001;
end_screen[38][30] = 16'b01011_011000_00100;
end_screen[38][31] = 16'b10100_100011_01010;
end_screen[38][32] = 16'b10111_100010_01001;
end_screen[38][33] = 16'b10011_011001_00100;
end_screen[38][34] = 16'b10001_010100_00010;
end_screen[38][35] = 16'b10000_010010_00010;
end_screen[38][36] = 16'b10000_010010_00010;
end_screen[38][37] = 16'b10000_010010_00010;
end_screen[38][38] = 16'b10000_010010_00010;
end_screen[38][39] = 16'b10100_101001_10100;
end_screen[38][40] = 16'b10100_101001_10100;
end_screen[38][41] = 16'b11111_111111_11111;
end_screen[38][42] = 16'b11111_111111_11111;
end_screen[38][43] = 16'b11111_111111_11111;
end_screen[38][44] = 16'b11111_111111_11111;
end_screen[38][45] = 16'b10100_101001_10100;
end_screen[38][46] = 16'b10100_101001_10100;
end_screen[38][47] = 16'b10100_101001_10100;
end_screen[38][48] = 16'b11111_111111_11111;
end_screen[38][49] = 16'b11111_111111_11111;
end_screen[38][50] = 16'b11111_111111_11111;
end_screen[38][51] = 16'b11111_111111_11111;
end_screen[38][52] = 16'b10100_101001_10100;
end_screen[38][53] = 16'b10100_101001_10100;
end_screen[38][54] = 16'b10100_101001_10100;
end_screen[38][55] = 16'b11111_111111_11111;
end_screen[38][56] = 16'b11111_111111_11111;
end_screen[38][57] = 16'b11111_111111_11111;
end_screen[38][58] = 16'b11001_010000_00001;
end_screen[38][59] = 16'b11001_010000_00001;
end_screen[38][60] = 16'b11010_010011_00010;
end_screen[38][61] = 16'b11010_010011_00010;
end_screen[38][62] = 16'b11010_010011_00010;
end_screen[38][63] = 16'b11010_010011_00010;
end_screen[38][64] = 16'b11001_010110_00100;
end_screen[38][65] = 16'b11010_100011_01010;
end_screen[38][66] = 16'b11010_101100_01111;
end_screen[38][67] = 16'b11001_101011_01101;
end_screen[38][68] = 16'b11001_101001_01101;
end_screen[38][69] = 16'b11001_100100_01011;
end_screen[38][70] = 16'b10111_010100_00100;
end_screen[38][71] = 16'b10110_000110_00000;
end_screen[38][72] = 16'b10111_000101_00000;
end_screen[38][73] = 16'b11000_001001_00000;
end_screen[38][74] = 16'b11000_001100_00001;
end_screen[38][75] = 16'b11000_001100_00001;
end_screen[38][76] = 16'b11000_001101_00001;
end_screen[38][77] = 16'b11000_001101_00001;
end_screen[38][78] = 16'b11001_001110_00001;
end_screen[38][79] = 16'b11001_001111_00010;
end_screen[38][80] = 16'b11001_001111_00010;
end_screen[38][81] = 16'b11001_001110_00001;
end_screen[38][82] = 16'b11010_001100_00001;
end_screen[38][83] = 16'b10101_010001_00010;
end_screen[38][84] = 16'b10010_010001_00001;
end_screen[38][85] = 16'b10111_001000_00000;
end_screen[38][86] = 16'b11010_000001_00000;
end_screen[38][87] = 16'b11000_000111_00000;
end_screen[38][88] = 16'b11000_010100_00011;
end_screen[38][89] = 16'b11001_100011_01010;
end_screen[38][90] = 16'b11001_101000_01100;
end_screen[38][91] = 16'b11001_101001_01101;
end_screen[38][92] = 16'b11010_101110_10000;
end_screen[38][93] = 16'b11000_101111_10101;
end_screen[38][94] = 16'b10011_101011_11011;
end_screen[38][95] = 16'b10001_101010_11100;
end_screen[39][0] = 16'b10001_101010_11100;
end_screen[39][1] = 16'b10001_101010_11100;
end_screen[39][2] = 16'b10001_101010_11100;
end_screen[39][3] = 16'b10011_101011_11011;
end_screen[39][4] = 16'b11001_101110_10010;
end_screen[39][5] = 16'b11101_110010_10001;
end_screen[39][6] = 16'b11100_110001_10001;
end_screen[39][7] = 16'b11010_101100_01110;
end_screen[39][8] = 16'b11010_100110_01000;
end_screen[39][9] = 16'b11011_100001_00010;
end_screen[39][10] = 16'b11100_100111_00111;
end_screen[39][11] = 16'b11101_101101_01011;
end_screen[39][12] = 16'b11100_100111_00110;
end_screen[39][13] = 16'b11010_100011_00101;
end_screen[39][14] = 16'b11001_011111_00100;
end_screen[39][15] = 16'b10111_011101_00100;
end_screen[39][16] = 16'b10111_011001_00000;
end_screen[39][17] = 16'b11000_011111_00100;
end_screen[39][18] = 16'b11100_110001_10010;
end_screen[39][19] = 16'b11111_111100_11000;
end_screen[39][20] = 16'b11110_111000_10110;
end_screen[39][21] = 16'b11110_111000_10110;
end_screen[39][22] = 16'b11110_110111_10110;
end_screen[39][23] = 16'b11101_110101_10100;
end_screen[39][24] = 16'b11101_110110_10101;
end_screen[39][25] = 16'b11111_111001_10111;
end_screen[39][26] = 16'b11111_111001_10110;
end_screen[39][27] = 16'b11110_110111_10101;
end_screen[39][28] = 16'b11011_110001_10001;
end_screen[39][29] = 16'b01111_100000_00111;
end_screen[39][30] = 16'b01001_010101_00010;
end_screen[39][31] = 16'b10100_100011_01010;
end_screen[39][32] = 16'b11100_101111_01111;
end_screen[39][33] = 16'b11001_100110_01011;
end_screen[39][34] = 16'b10001_010101_00011;
end_screen[39][35] = 16'b10001_010100_00011;
end_screen[39][36] = 16'b10001_010101_00011;
end_screen[39][37] = 16'b10001_010100_00011;
end_screen[39][38] = 16'b10001_010100_00011;
end_screen[39][39] = 16'b10100_101001_10100;
end_screen[39][40] = 16'b10100_101001_10100;
end_screen[39][41] = 16'b11111_111111_11111;
end_screen[39][42] = 16'b11111_111111_11111;
end_screen[39][43] = 16'b11111_111111_11111;
end_screen[39][44] = 16'b11111_111111_11111;
end_screen[39][45] = 16'b10100_101001_10100;
end_screen[39][46] = 16'b10100_101001_10100;
end_screen[39][47] = 16'b10100_101001_10100;
end_screen[39][48] = 16'b11111_111111_11111;
end_screen[39][49] = 16'b11111_111111_11111;
end_screen[39][50] = 16'b11111_111111_11111;
end_screen[39][51] = 16'b11111_111111_11111;
end_screen[39][52] = 16'b10100_101001_10100;
end_screen[39][53] = 16'b10100_101001_10100;
end_screen[39][54] = 16'b10100_101001_10100;
end_screen[39][55] = 16'b11111_111111_11111;
end_screen[39][56] = 16'b11111_111111_11111;
end_screen[39][57] = 16'b11111_111111_11111;
end_screen[39][58] = 16'b11001_010111_00100;
end_screen[39][59] = 16'b11001_010111_00100;
end_screen[39][60] = 16'b11001_010011_00010;
end_screen[39][61] = 16'b11000_001101_00000;
end_screen[39][62] = 16'b10111_001010_00000;
end_screen[39][63] = 16'b11000_001110_00000;
end_screen[39][64] = 16'b11010_100000_01001;
end_screen[39][65] = 16'b11001_101010_01101;
end_screen[39][66] = 16'b11001_101011_01110;
end_screen[39][67] = 16'b11001_101000_01100;
end_screen[39][68] = 16'b11000_011100_00111;
end_screen[39][69] = 16'b10111_001001_00000;
end_screen[39][70] = 16'b10110_000111_00000;
end_screen[39][71] = 16'b10111_001011_00001;
end_screen[39][72] = 16'b11000_001101_00001;
end_screen[39][73] = 16'b11010_010000_00010;
end_screen[39][74] = 16'b11001_010000_00010;
end_screen[39][75] = 16'b11001_001110_00001;
end_screen[39][76] = 16'b11000_001110_00001;
end_screen[39][77] = 16'b11001_001110_00001;
end_screen[39][78] = 16'b11001_001110_00001;
end_screen[39][79] = 16'b11001_001111_00010;
end_screen[39][80] = 16'b11001_001110_00001;
end_screen[39][81] = 16'b11001_001110_00001;
end_screen[39][82] = 16'b10101_010001_00010;
end_screen[39][83] = 16'b01011_011011_00011;
end_screen[39][84] = 16'b01000_011110_00011;
end_screen[39][85] = 16'b10000_010010_00001;
end_screen[39][86] = 16'b10100_001011_00000;
end_screen[39][87] = 16'b10101_001010_00000;
end_screen[39][88] = 16'b11000_000111_00000;
end_screen[39][89] = 16'b10111_001010_00000;
end_screen[39][90] = 16'b11000_011010_00110;
end_screen[39][91] = 16'b11001_101000_01100;
end_screen[39][92] = 16'b11010_101110_10000;
end_screen[39][93] = 16'b11011_110000_10001;
end_screen[39][94] = 16'b10111_101111_10111;
end_screen[39][95] = 16'b10001_101010_11100;
end_screen[40][0] = 16'b10001_101010_11100;
end_screen[40][1] = 16'b10001_101010_11100;
end_screen[40][2] = 16'b10100_101101_11001;
end_screen[40][3] = 16'b11010_110000_10011;
end_screen[40][4] = 16'b11100_101111_01111;
end_screen[40][5] = 16'b11100_110010_10010;
end_screen[40][6] = 16'b11100_110010_10010;
end_screen[40][7] = 16'b11010_100101_00111;
end_screen[40][8] = 16'b11011_011111_00001;
end_screen[40][9] = 16'b11011_100010_00011;
end_screen[40][10] = 16'b11011_100101_00110;
end_screen[40][11] = 16'b11011_100011_00100;
end_screen[40][12] = 16'b11010_011111_00001;
end_screen[40][13] = 16'b11010_100001_00011;
end_screen[40][14] = 16'b11001_011110_00010;
end_screen[40][15] = 16'b11000_011100_00001;
end_screen[40][16] = 16'b11000_011001_00000;
end_screen[40][17] = 16'b11000_011011_00010;
end_screen[40][18] = 16'b11011_101010_01100;
end_screen[40][19] = 16'b11110_111001_10111;
end_screen[40][20] = 16'b11110_110111_10110;
end_screen[40][21] = 16'b11101_110110_10100;
end_screen[40][22] = 16'b11110_110111_10101;
end_screen[40][23] = 16'b11110_110111_10101;
end_screen[40][24] = 16'b11101_110110_10100;
end_screen[40][25] = 16'b11101_110110_10100;
end_screen[40][26] = 16'b11101_110110_10101;
end_screen[40][27] = 16'b11110_110110_10100;
end_screen[40][28] = 16'b11110_110101_10100;
end_screen[40][29] = 16'b11000_101101_01111;
end_screen[40][30] = 16'b01101_011101_00110;
end_screen[40][31] = 16'b10100_100100_01010;
end_screen[40][32] = 16'b11100_101110_01111;
end_screen[40][33] = 16'b11100_101111_10000;
end_screen[40][34] = 16'b11000_100110_01011;
end_screen[40][35] = 16'b10101_011101_00110;
end_screen[40][36] = 16'b10110_011110_00110;
end_screen[40][37] = 16'b10110_011101_00110;
end_screen[40][38] = 16'b10110_011101_00110;
end_screen[40][39] = 16'b11111_110011_00111;
end_screen[40][40] = 16'b11111_110011_00111;
end_screen[40][41] = 16'b11111_110011_00111;
end_screen[40][42] = 16'b11111_110011_00111;
end_screen[40][43] = 16'b11111_110011_00111;
end_screen[40][44] = 16'b11111_110011_00111;
end_screen[40][45] = 16'b11111_110011_00111;
end_screen[40][46] = 16'b11111_110011_00111;
end_screen[40][47] = 16'b11111_110011_00111;
end_screen[40][48] = 16'b11111_110011_00111;
end_screen[40][49] = 16'b11111_110011_00111;
end_screen[40][50] = 16'b11111_110011_00111;
end_screen[40][51] = 16'b11111_110011_00111;
end_screen[40][52] = 16'b11111_110011_00111;
end_screen[40][53] = 16'b11111_110011_00111;
end_screen[40][54] = 16'b11111_110011_00111;
end_screen[40][55] = 16'b11111_110011_00111;
end_screen[40][56] = 16'b11111_110011_00111;
end_screen[40][57] = 16'b11111_110011_00111;
end_screen[40][58] = 16'b11001_100100_01010;
end_screen[40][59] = 16'b11001_100100_01010;
end_screen[40][60] = 16'b11001_100001_01000;
end_screen[40][61] = 16'b11001_011110_01000;
end_screen[40][62] = 16'b11000_011011_00110;
end_screen[40][63] = 16'b11000_011101_00111;
end_screen[40][64] = 16'b11010_100110_01100;
end_screen[40][65] = 16'b11010_101101_01111;
end_screen[40][66] = 16'b11001_100111_01100;
end_screen[40][67] = 16'b11000_011000_00101;
end_screen[40][68] = 16'b10111_001010_00000;
end_screen[40][69] = 16'b10110_001001_00000;
end_screen[40][70] = 16'b11000_001101_00001;
end_screen[40][71] = 16'b11001_001111_00010;
end_screen[40][72] = 16'b11001_001111_00010;
end_screen[40][73] = 16'b11001_001111_00001;
end_screen[40][74] = 16'b11000_001101_00001;
end_screen[40][75] = 16'b11000_001101_00001;
end_screen[40][76] = 16'b11000_001101_00001;
end_screen[40][77] = 16'b11000_001101_00001;
end_screen[40][78] = 16'b11000_001101_00001;
end_screen[40][79] = 16'b11000_001101_00001;
end_screen[40][80] = 16'b11001_001011_00001;
end_screen[40][81] = 16'b10101_001111_00001;
end_screen[40][82] = 16'b01001_011100_00011;
end_screen[40][83] = 16'b01011_011011_00011;
end_screen[40][84] = 16'b01011_011001_00011;
end_screen[40][85] = 16'b01010_011000_00010;
end_screen[40][86] = 16'b00110_011001_00010;
end_screen[40][87] = 16'b01110_010010_00001;
end_screen[40][88] = 16'b11000_001010_00001;
end_screen[40][89] = 16'b10111_001010_00000;
end_screen[40][90] = 16'b10111_001010_00000;
end_screen[40][91] = 16'b11000_011001_00101;
end_screen[40][92] = 16'b11001_101001_01100;
end_screen[40][93] = 16'b11011_110001_10010;
end_screen[40][94] = 16'b10111_110000_11000;
end_screen[40][95] = 16'b10001_101010_11100;
end_screen[41][0] = 16'b10001_101010_11100;
end_screen[41][1] = 16'b10001_101010_11100;
end_screen[41][2] = 16'b10111_101111_10110;
end_screen[41][3] = 16'b11100_110001_10000;
end_screen[41][4] = 16'b11100_110010_10010;
end_screen[41][5] = 16'b11100_110001_10000;
end_screen[41][6] = 16'b11100_101011_01010;
end_screen[41][7] = 16'b11010_100000_00010;
end_screen[41][8] = 16'b11001_011101_00000;
end_screen[41][9] = 16'b11010_100000_00011;
end_screen[41][10] = 16'b11010_100001_00011;
end_screen[41][11] = 16'b11010_100010_00100;
end_screen[41][12] = 16'b11011_100110_00111;
end_screen[41][13] = 16'b11100_101010_01000;
end_screen[41][14] = 16'b11100_101001_01000;
end_screen[41][15] = 16'b11011_100101_00101;
end_screen[41][16] = 16'b11010_100011_00100;
end_screen[41][17] = 16'b11001_011011_00000;
end_screen[41][18] = 16'b11010_011111_00010;
end_screen[41][19] = 16'b11100_101111_01111;
end_screen[41][20] = 16'b11101_110110_10100;
end_screen[41][21] = 16'b11101_110100_10011;
end_screen[41][22] = 16'b11110_110111_10101;
end_screen[41][23] = 16'b11110_110111_10101;
end_screen[41][24] = 16'b11101_110011_10011;
end_screen[41][25] = 16'b11101_110100_10011;
end_screen[41][26] = 16'b11101_110110_10100;
end_screen[41][27] = 16'b11101_110101_10011;
end_screen[41][28] = 16'b11101_110101_10100;
end_screen[41][29] = 16'b11111_110111_10101;
end_screen[41][30] = 16'b11000_101100_01110;
end_screen[41][31] = 16'b11000_101010_01101;
end_screen[41][32] = 16'b11100_101111_10000;
end_screen[41][33] = 16'b11011_101110_01111;
end_screen[41][34] = 16'b11010_101100_01110;
end_screen[41][35] = 16'b10101_011011_00101;
end_screen[41][36] = 16'b10101_011101_00110;
end_screen[41][37] = 16'b10110_011110_00110;
end_screen[41][38] = 16'b10110_011110_00110;
end_screen[41][39] = 16'b11111_110011_00111;
end_screen[41][40] = 16'b11111_110011_00111;
end_screen[41][41] = 16'b11111_110011_00111;
end_screen[41][42] = 16'b11111_110011_00111;
end_screen[41][43] = 16'b11111_110011_00111;
end_screen[41][44] = 16'b11111_110011_00111;
end_screen[41][45] = 16'b11111_110011_00111;
end_screen[41][46] = 16'b11111_110011_00111;
end_screen[41][47] = 16'b11111_110011_00111;
end_screen[41][48] = 16'b11111_110011_00111;
end_screen[41][49] = 16'b11111_110011_00111;
end_screen[41][50] = 16'b11111_110011_00111;
end_screen[41][51] = 16'b11111_110011_00111;
end_screen[41][52] = 16'b11111_110011_00111;
end_screen[41][53] = 16'b11111_110011_00111;
end_screen[41][54] = 16'b11111_110011_00111;
end_screen[41][55] = 16'b11111_110011_00111;
end_screen[41][56] = 16'b11111_110011_00111;
end_screen[41][57] = 16'b11111_110011_00111;
end_screen[41][58] = 16'b11010_101101_01110;
end_screen[41][59] = 16'b11010_101101_01110;
end_screen[41][60] = 16'b11010_101110_01111;
end_screen[41][61] = 16'b11010_110000_10000;
end_screen[41][62] = 16'b11010_101111_01111;
end_screen[41][63] = 16'b11011_110010_10011;
end_screen[41][64] = 16'b11011_110001_10010;
end_screen[41][65] = 16'b11001_101000_01100;
end_screen[41][66] = 16'b11000_011011_00110;
end_screen[41][67] = 16'b10111_001011_00000;
end_screen[41][68] = 16'b10111_001010_00000;
end_screen[41][69] = 16'b10111_001011_00001;
end_screen[41][70] = 16'b11000_001110_00001;
end_screen[41][71] = 16'b11010_010000_00010;
end_screen[41][72] = 16'b11001_001111_00010;
end_screen[41][73] = 16'b11001_001110_00001;
end_screen[41][74] = 16'b11000_001101_00001;
end_screen[41][75] = 16'b11000_001101_00001;
end_screen[41][76] = 16'b11000_001101_00001;
end_screen[41][77] = 16'b11000_001101_00001;
end_screen[41][78] = 16'b11000_001101_00001;
end_screen[41][79] = 16'b11000_001110_00001;
end_screen[41][80] = 16'b11001_001011_00001;
end_screen[41][81] = 16'b10101_001110_00001;
end_screen[41][82] = 16'b01011_011010_00011;
end_screen[41][83] = 16'b01011_011011_00011;
end_screen[41][84] = 16'b01011_011001_00011;
end_screen[41][85] = 16'b01100_011100_00011;
end_screen[41][86] = 16'b01101_011110_00100;
end_screen[41][87] = 16'b01011_011110_00011;
end_screen[41][88] = 16'b01110_010110_00010;
end_screen[41][89] = 16'b11000_001010_00001;
end_screen[41][90] = 16'b11000_001100_00001;
end_screen[41][91] = 16'b10111_001000_00000;
end_screen[41][92] = 16'b11000_011110_01000;
end_screen[41][93] = 16'b11011_110001_10010;
end_screen[41][94] = 16'b10111_110000_11001;
end_screen[41][95] = 16'b10001_101010_11100;
end_screen[42][0] = 16'b10001_101010_11100;
end_screen[42][1] = 16'b10100_101101_11010;
end_screen[42][2] = 16'b11001_110001_10101;
end_screen[42][3] = 16'b11100_110010_10001;
end_screen[42][4] = 16'b11100_110011_10010;
end_screen[42][5] = 16'b11011_101100_01101;
end_screen[42][6] = 16'b11001_011100_00000;
end_screen[42][7] = 16'b11001_011011_00000;
end_screen[42][8] = 16'b11001_011111_00011;
end_screen[42][9] = 16'b11010_100010_00100;
end_screen[42][10] = 16'b11100_101000_01000;
end_screen[42][11] = 16'b11101_101110_01100;
end_screen[42][12] = 16'b11101_101110_01100;
end_screen[42][13] = 16'b11100_101001_01001;
end_screen[42][14] = 16'b11100_101000_01000;
end_screen[42][15] = 16'b11010_100010_00100;
end_screen[42][16] = 16'b11001_011111_00010;
end_screen[42][17] = 16'b11001_011101_00010;
end_screen[42][18] = 16'b11000_011010_00000;
end_screen[42][19] = 16'b11010_100010_00100;
end_screen[42][20] = 16'b11101_110101_10100;
end_screen[42][21] = 16'b11101_110110_10101;
end_screen[42][22] = 16'b11101_110101_10100;
end_screen[42][23] = 16'b11101_110100_10011;
end_screen[42][24] = 16'b11101_110100_10011;
end_screen[42][25] = 16'b11101_110110_10101;
end_screen[42][26] = 16'b11110_110111_10101;
end_screen[42][27] = 16'b11101_110110_10100;
end_screen[42][28] = 16'b11101_110101_10100;
end_screen[42][29] = 16'b11101_110101_10011;
end_screen[42][30] = 16'b11110_110101_10011;
end_screen[42][31] = 16'b11011_101110_01111;
end_screen[42][32] = 16'b11010_101011_01110;
end_screen[42][33] = 16'b11011_101111_10000;
end_screen[42][34] = 16'b11010_101100_01110;
end_screen[42][35] = 16'b10110_100010_01001;
end_screen[42][36] = 16'b10101_011100_00101;
end_screen[42][37] = 16'b10100_011011_00101;
end_screen[42][38] = 16'b10100_011011_00101;
end_screen[42][39] = 16'b11111_110011_00111;
end_screen[42][40] = 16'b11111_110011_00111;
end_screen[42][41] = 16'b11111_110011_00111;
end_screen[42][42] = 16'b11111_110011_00111;
end_screen[42][43] = 16'b11111_110011_00111;
end_screen[42][44] = 16'b11111_110011_00111;
end_screen[42][45] = 16'b11111_110011_00111;
end_screen[42][46] = 16'b11111_110011_00111;
end_screen[42][47] = 16'b11111_110011_00111;
end_screen[42][48] = 16'b11111_110011_00111;
end_screen[42][49] = 16'b11111_110011_00111;
end_screen[42][50] = 16'b11111_110011_00111;
end_screen[42][51] = 16'b11111_110011_00111;
end_screen[42][52] = 16'b11111_110011_00111;
end_screen[42][53] = 16'b11111_110011_00111;
end_screen[42][54] = 16'b11111_110011_00111;
end_screen[42][55] = 16'b11111_110011_00111;
end_screen[42][56] = 16'b11111_110011_00111;
end_screen[42][57] = 16'b11111_110011_00111;
end_screen[42][58] = 16'b11100_110001_10001;
end_screen[42][59] = 16'b11100_110001_10001;
end_screen[42][60] = 16'b11100_110001_10001;
end_screen[42][61] = 16'b11011_101111_10000;
end_screen[42][62] = 16'b11011_101111_10000;
end_screen[42][63] = 16'b11100_110010_10011;
end_screen[42][64] = 16'b11011_110011_10011;
end_screen[42][65] = 16'b11001_100010_01010;
end_screen[42][66] = 16'b10111_001100_00000;
end_screen[42][67] = 16'b10111_001010_00000;
end_screen[42][68] = 16'b10111_001011_00001;
end_screen[42][69] = 16'b10111_001011_00001;
end_screen[42][70] = 16'b11001_001110_00001;
end_screen[42][71] = 16'b11010_010000_00010;
end_screen[42][72] = 16'b11001_001111_00010;
end_screen[42][73] = 16'b11000_001101_00001;
end_screen[42][74] = 16'b11000_001101_00001;
end_screen[42][75] = 16'b11001_001110_00001;
end_screen[42][76] = 16'b11001_001110_00001;
end_screen[42][77] = 16'b11000_001110_00001;
end_screen[42][78] = 16'b11001_001110_00001;
end_screen[42][79] = 16'b11001_001111_00010;
end_screen[42][80] = 16'b11001_001110_00001;
end_screen[42][81] = 16'b11001_001101_00001;
end_screen[42][82] = 16'b10110_001111_00001;
end_screen[42][83] = 16'b01011_011010_00011;
end_screen[42][84] = 16'b01010_011011_00011;
end_screen[42][85] = 16'b01011_011010_00011;
end_screen[42][86] = 16'b01100_011010_00011;
end_screen[42][87] = 16'b01001_011100_00011;
end_screen[42][88] = 16'b01011_010110_00010;
end_screen[42][89] = 16'b11001_001011_00001;
end_screen[42][90] = 16'b11001_001111_00010;
end_screen[42][91] = 16'b10111_001001_00000;
end_screen[42][92] = 16'b10110_001110_00001;
end_screen[42][93] = 16'b11010_100111_01101;
end_screen[42][94] = 16'b10111_110001_11001;
end_screen[42][95] = 16'b10001_101010_11100;
end_screen[43][0] = 16'b10001_101010_11100;
end_screen[43][1] = 16'b11010_110000_10011;
end_screen[43][2] = 16'b11101_110011_10010;
end_screen[43][3] = 16'b11101_110011_10010;
end_screen[43][4] = 16'b11011_101110_01111;
end_screen[43][5] = 16'b11001_100010_00111;
end_screen[43][6] = 16'b11000_011000_00000;
end_screen[43][7] = 16'b11001_011101_00010;
end_screen[43][8] = 16'b11100_100111_00111;
end_screen[43][9] = 16'b11101_101011_01001;
end_screen[43][10] = 16'b11101_101011_01001;
end_screen[43][11] = 16'b11100_101010_01001;
end_screen[43][12] = 16'b11011_100110_00110;
end_screen[43][13] = 16'b11010_100000_00011;
end_screen[43][14] = 16'b11001_011101_00001;
end_screen[43][15] = 16'b11010_011111_00011;
end_screen[43][16] = 16'b11000_011101_00010;
end_screen[43][17] = 16'b10111_011001_00000;
end_screen[43][18] = 16'b10111_010101_00000;
end_screen[43][19] = 16'b11000_011011_00001;
end_screen[43][20] = 16'b11101_110001_10001;
end_screen[43][21] = 16'b11110_110111_10101;
end_screen[43][22] = 16'b11101_110101_10100;
end_screen[43][23] = 16'b11101_110100_10011;
end_screen[43][24] = 16'b11110_110110_10101;
end_screen[43][25] = 16'b11110_110111_10101;
end_screen[43][26] = 16'b11101_110101_10100;
end_screen[43][27] = 16'b11101_110011_10010;
end_screen[43][28] = 16'b11101_110100_10011;
end_screen[43][29] = 16'b11101_110100_10011;
end_screen[43][30] = 16'b11101_110101_10100;
end_screen[43][31] = 16'b11011_101110_01111;
end_screen[43][32] = 16'b11010_101001_01100;
end_screen[43][33] = 16'b11011_101110_01111;
end_screen[43][34] = 16'b11100_110001_10001;
end_screen[43][35] = 16'b11100_110000_10001;
end_screen[43][36] = 16'b10001_010101_00011;
end_screen[43][37] = 16'b10001_010100_00010;
end_screen[43][38] = 16'b10001_010100_00010;
end_screen[43][39] = 16'b11111_110011_00111;
end_screen[43][40] = 16'b11111_110011_00111;
end_screen[43][41] = 16'b11111_110011_00111;
end_screen[43][42] = 16'b00000_000000_00000;
end_screen[43][43] = 16'b00000_000000_00000;
end_screen[43][44] = 16'b00000_000000_00000;
end_screen[43][45] = 16'b11111_110011_00111;
end_screen[43][46] = 16'b11111_110011_00111;
end_screen[43][47] = 16'b11111_110011_00111;
end_screen[43][48] = 16'b11111_110011_00111;
end_screen[43][49] = 16'b11111_110011_00111;
end_screen[43][50] = 16'b11111_110011_00111;
end_screen[43][51] = 16'b11111_110011_00111;
end_screen[43][52] = 16'b00000_000000_00000;
end_screen[43][53] = 16'b00000_000000_00000;
end_screen[43][54] = 16'b00000_000000_00000;
end_screen[43][55] = 16'b11111_110011_00111;
end_screen[43][56] = 16'b11111_110011_00111;
end_screen[43][57] = 16'b11111_110011_00111;
end_screen[43][58] = 16'b11011_101110_01111;
end_screen[43][59] = 16'b11011_101110_01111;
end_screen[43][60] = 16'b11011_101101_01111;
end_screen[43][61] = 16'b11010_101101_01111;
end_screen[43][62] = 16'b11011_101101_01111;
end_screen[43][63] = 16'b11011_110001_10010;
end_screen[43][64] = 16'b11100_110101_10100;
end_screen[43][65] = 16'b11001_100011_01100;
end_screen[43][66] = 16'b10110_000110_00000;
end_screen[43][67] = 16'b10111_001011_00000;
end_screen[43][68] = 16'b10111_001011_00001;
end_screen[43][69] = 16'b11000_001110_00001;
end_screen[43][70] = 16'b11001_001111_00010;
end_screen[43][71] = 16'b11001_010000_00010;
end_screen[43][72] = 16'b11001_001110_00001;
end_screen[43][73] = 16'b11000_001101_00001;
end_screen[43][74] = 16'b11000_001101_00001;
end_screen[43][75] = 16'b11001_001111_00010;
end_screen[43][76] = 16'b11001_001111_00010;
end_screen[43][77] = 16'b11001_001111_00001;
end_screen[43][78] = 16'b11001_001111_00010;
end_screen[43][79] = 16'b11001_001111_00010;
end_screen[43][80] = 16'b11001_001111_00001;
end_screen[43][81] = 16'b11010_001111_00010;
end_screen[43][82] = 16'b11010_001110_00001;
end_screen[43][83] = 16'b10110_001111_00001;
end_screen[43][84] = 16'b10110_001101_00001;
end_screen[43][85] = 16'b01110_010110_00010;
end_screen[43][86] = 16'b00111_100001_00100;
end_screen[43][87] = 16'b01110_010101_00010;
end_screen[43][88] = 16'b10111_001011_00000;
end_screen[43][89] = 16'b11000_001101_00001;
end_screen[43][90] = 16'b11001_001111_00010;
end_screen[43][91] = 16'b10111_001011_00001;
end_screen[43][92] = 16'b10110_000111_00000;
end_screen[43][93] = 16'b11001_100010_01011;
end_screen[43][94] = 16'b10111_110001_11001;
end_screen[43][95] = 16'b10001_101010_11100;
end_screen[44][0] = 16'b10001_101010_11100;
end_screen[44][1] = 16'b11001_110000_10101;
end_screen[44][2] = 16'b11101_110011_10010;
end_screen[44][3] = 16'b11100_110011_10011;
end_screen[44][4] = 16'b11001_100110_01010;
end_screen[44][5] = 16'b10111_010111_00000;
end_screen[44][6] = 16'b11011_100000_00010;
end_screen[44][7] = 16'b11100_101000_00111;
end_screen[44][8] = 16'b11100_101001_01000;
end_screen[44][9] = 16'b11100_100111_00111;
end_screen[44][10] = 16'b11011_100011_00011;
end_screen[44][11] = 16'b11010_011101_00000;
end_screen[44][12] = 16'b11010_011101_00001;
end_screen[44][13] = 16'b11010_100001_00100;
end_screen[44][14] = 16'b11011_100100_00110;
end_screen[44][15] = 16'b11011_100110_00111;
end_screen[44][16] = 16'b11011_101000_01000;
end_screen[44][17] = 16'b11010_100010_00100;
end_screen[44][18] = 16'b10111_010111_00000;
end_screen[44][19] = 16'b10111_010111_00000;
end_screen[44][20] = 16'b11100_101000_00111;
end_screen[44][21] = 16'b11101_110101_10011;
end_screen[44][22] = 16'b11110_110111_10110;
end_screen[44][23] = 16'b11101_110101_10100;
end_screen[44][24] = 16'b11101_110101_10100;
end_screen[44][25] = 16'b11101_110101_10100;
end_screen[44][26] = 16'b11100_110011_10010;
end_screen[44][27] = 16'b11101_110100_10011;
end_screen[44][28] = 16'b11101_110110_10100;
end_screen[44][29] = 16'b11101_110110_10100;
end_screen[44][30] = 16'b11101_110100_10011;
end_screen[44][31] = 16'b11100_110010_10010;
end_screen[44][32] = 16'b11010_101010_01101;
end_screen[44][33] = 16'b11010_101001_01100;
end_screen[44][34] = 16'b11100_110010_10001;
end_screen[44][35] = 16'b11011_110001_10001;
end_screen[44][36] = 16'b10001_100101_10101;
end_screen[44][37] = 16'b10001_100101_10101;
end_screen[44][38] = 16'b10001_101010_11100;
end_screen[44][39] = 16'b11111_110011_00111;
end_screen[44][40] = 16'b11111_110011_00111;
end_screen[44][41] = 16'b11111_110011_00111;
end_screen[44][42] = 16'b00000_000000_00000;
end_screen[44][43] = 16'b00000_000000_00000;
end_screen[44][44] = 16'b00000_000000_00000;
end_screen[44][45] = 16'b11111_110011_00111;
end_screen[44][46] = 16'b11111_110011_00111;
end_screen[44][47] = 16'b11111_110011_00111;
end_screen[44][48] = 16'b11111_110011_00111;
end_screen[44][49] = 16'b11111_110011_00111;
end_screen[44][50] = 16'b11111_110011_00111;
end_screen[44][51] = 16'b11111_110011_00111;
end_screen[44][52] = 16'b00000_000000_00000;
end_screen[44][53] = 16'b00000_000000_00000;
end_screen[44][54] = 16'b00000_000000_00000;
end_screen[44][55] = 16'b11111_110011_00111;
end_screen[44][56] = 16'b11111_110100_01000;
end_screen[44][57] = 16'b11111_110011_00111;
end_screen[44][58] = 16'b10101_100111_10010;
end_screen[44][59] = 16'b10101_100111_10010;
end_screen[44][60] = 16'b10101_101001_10010;
end_screen[44][61] = 16'b10110_101010_10011;
end_screen[44][62] = 16'b10110_101001_10011;
end_screen[44][63] = 16'b11001_101110_10011;
end_screen[44][64] = 16'b11100_111000_10110;
end_screen[44][65] = 16'b11010_100101_01110;
end_screen[44][66] = 16'b10110_000011_00000;
end_screen[44][67] = 16'b10111_001011_00000;
end_screen[44][68] = 16'b10111_001100_00001;
end_screen[44][69] = 16'b11001_001110_00001;
end_screen[44][70] = 16'b11001_001111_00010;
end_screen[44][71] = 16'b11001_001111_00010;
end_screen[44][72] = 16'b11001_001111_00010;
end_screen[44][73] = 16'b11000_001100_00001;
end_screen[44][74] = 16'b11000_001100_00001;
end_screen[44][75] = 16'b11001_001110_00001;
end_screen[44][76] = 16'b11001_001110_00001;
end_screen[44][77] = 16'b11001_001110_00001;
end_screen[44][78] = 16'b11000_001101_00001;
end_screen[44][79] = 16'b11001_001110_00001;
end_screen[44][80] = 16'b11001_001111_00010;
end_screen[44][81] = 16'b11001_001111_00010;
end_screen[44][82] = 16'b11001_001111_00010;
end_screen[44][83] = 16'b11001_001100_00001;
end_screen[44][84] = 16'b11010_001001_00000;
end_screen[44][85] = 16'b10101_001110_00001;
end_screen[44][86] = 16'b10001_010011_00010;
end_screen[44][87] = 16'b10110_001110_00001;
end_screen[44][88] = 16'b11010_001011_00001;
end_screen[44][89] = 16'b11000_001110_00001;
end_screen[44][90] = 16'b11001_001111_00010;
end_screen[44][91] = 16'b10111_000111_00000;
end_screen[44][92] = 16'b10111_010011_00011;
end_screen[44][93] = 16'b11010_101010_01110;
end_screen[44][94] = 16'b10111_101111_11000;
end_screen[44][95] = 16'b10001_101010_11100;
end_screen[45][0] = 16'b10001_101010_11100;
end_screen[45][1] = 16'b11001_110001_10101;
end_screen[45][2] = 16'b11101_110011_10010;
end_screen[45][3] = 16'b11100_110010_10010;
end_screen[45][4] = 16'b11001_100100_01001;
end_screen[45][5] = 16'b10111_011000_00000;
end_screen[45][6] = 16'b11011_100000_00010;
end_screen[45][7] = 16'b11100_100100_00100;
end_screen[45][8] = 16'b11011_100001_00010;
end_screen[45][9] = 16'b11001_011011_00000;
end_screen[45][10] = 16'b11010_011011_00000;
end_screen[45][11] = 16'b11011_100011_00011;
end_screen[45][12] = 16'b11101_101100_01010;
end_screen[45][13] = 16'b11101_110001_10000;
end_screen[45][14] = 16'b11101_110001_10000;
end_screen[45][15] = 16'b11100_101011_01010;
end_screen[45][16] = 16'b11100_101000_01000;
end_screen[45][17] = 16'b11010_100010_00100;
end_screen[45][18] = 16'b11000_011010_00000;
end_screen[45][19] = 16'b11001_011011_00000;
end_screen[45][20] = 16'b11100_101000_01000;
end_screen[45][21] = 16'b11101_110011_10010;
end_screen[45][22] = 16'b11101_110101_10100;
end_screen[45][23] = 16'b11110_110110_10101;
end_screen[45][24] = 16'b11101_110100_10011;
end_screen[45][25] = 16'b11100_110010_10010;
end_screen[45][26] = 16'b11101_110100_10011;
end_screen[45][27] = 16'b11110_110110_10100;
end_screen[45][28] = 16'b11101_110100_10011;
end_screen[45][29] = 16'b11101_110011_10010;
end_screen[45][30] = 16'b11101_110100_10011;
end_screen[45][31] = 16'b11101_110100_10011;
end_screen[45][32] = 16'b11010_101011_01101;
end_screen[45][33] = 16'b11001_101001_01100;
end_screen[45][34] = 16'b11100_110010_10001;
end_screen[45][35] = 16'b11011_110001_10010;
end_screen[45][36] = 16'b10001_101010_11100;
end_screen[45][37] = 16'b10001_101010_11100;
end_screen[45][38] = 16'b10001_101010_11100;
end_screen[45][39] = 16'b11111_110011_00111;
end_screen[45][40] = 16'b11111_110011_00111;
end_screen[45][41] = 16'b11111_110011_00111;
end_screen[45][42] = 16'b00000_000000_00000;
end_screen[45][43] = 16'b00000_000000_00000;
end_screen[45][44] = 16'b00000_000000_00000;
end_screen[45][45] = 16'b11111_110011_00111;
end_screen[45][46] = 16'b11111_110011_00111;
end_screen[45][47] = 16'b11111_110011_00111;
end_screen[45][48] = 16'b11111_110011_00111;
end_screen[45][49] = 16'b11111_110011_00111;
end_screen[45][50] = 16'b11111_110011_00111;
end_screen[45][51] = 16'b11111_110011_00111;
end_screen[45][52] = 16'b00000_000000_00000;
end_screen[45][53] = 16'b00000_000000_00000;
end_screen[45][54] = 16'b00000_000000_00000;
end_screen[45][55] = 16'b11111_110011_00111;
end_screen[45][56] = 16'b11111_110100_01000;
end_screen[45][57] = 16'b11111_110011_00111;
end_screen[45][58] = 16'b10001_101010_11100;
end_screen[45][59] = 16'b10001_101010_11100;
end_screen[45][60] = 16'b10001_101010_11100;
end_screen[45][61] = 16'b10001_101010_11100;
end_screen[45][62] = 16'b10001_101010_11100;
end_screen[45][63] = 16'b11000_101110_10101;
end_screen[45][64] = 16'b11100_110011_10100;
end_screen[45][65] = 16'b11011_101011_01111;
end_screen[45][66] = 16'b10111_010000_00010;
end_screen[45][67] = 16'b10111_000111_00000;
end_screen[45][68] = 16'b10111_001010_00000;
end_screen[45][69] = 16'b10111_001100_00001;
end_screen[45][70] = 16'b11001_001111_00001;
end_screen[45][71] = 16'b11010_010000_00010;
end_screen[45][72] = 16'b11001_001111_00010;
end_screen[45][73] = 16'b11000_001101_00001;
end_screen[45][74] = 16'b11000_001101_00001;
end_screen[45][75] = 16'b11000_001101_00001;
end_screen[45][76] = 16'b11000_001110_00001;
end_screen[45][77] = 16'b11000_001110_00001;
end_screen[45][78] = 16'b11000_001101_00001;
end_screen[45][79] = 16'b11000_001100_00001;
end_screen[45][80] = 16'b11000_001101_00001;
end_screen[45][81] = 16'b11000_001101_00001;
end_screen[45][82] = 16'b10111_001100_00001;
end_screen[45][83] = 16'b10111_001011_00001;
end_screen[45][84] = 16'b10111_001011_00001;
end_screen[45][85] = 16'b11000_001001_00000;
end_screen[45][86] = 16'b11010_001000_00000;
end_screen[45][87] = 16'b11010_001101_00001;
end_screen[45][88] = 16'b11001_010000_00010;
end_screen[45][89] = 16'b11001_001101_00001;
end_screen[45][90] = 16'b11000_001001_00000;
end_screen[45][91] = 16'b10110_001011_00000;
end_screen[45][92] = 16'b11010_101000_01110;
end_screen[45][93] = 16'b11011_110001_10010;
end_screen[45][94] = 16'b10110_101011_10101;
end_screen[45][95] = 16'b10001_101010_11100;
end_screen[46][0] = 16'b10001_101010_11100;
end_screen[46][1] = 16'b11001_110000_10101;
end_screen[46][2] = 16'b11101_110100_10011;
end_screen[46][3] = 16'b11100_110011_10010;
end_screen[46][4] = 16'b11001_100100_01010;
end_screen[46][5] = 16'b10111_010111_00000;
end_screen[46][6] = 16'b11011_100000_00001;
end_screen[46][7] = 16'b10111_011000_00000;
end_screen[46][8] = 16'b10101_010011_00000;
end_screen[46][9] = 16'b11001_011100_00000;
end_screen[46][10] = 16'b11101_100111_00101;
end_screen[46][11] = 16'b11101_101101_01010;
end_screen[46][12] = 16'b11110_101111_01100;
end_screen[46][13] = 16'b11101_101100_01001;
end_screen[46][14] = 16'b11100_101010_01001;
end_screen[46][15] = 16'b11010_100100_00110;
end_screen[46][16] = 16'b11010_100011_00110;
end_screen[46][17] = 16'b11001_100000_00100;
end_screen[46][18] = 16'b10111_011001_00001;
end_screen[46][19] = 16'b11000_011011_00001;
end_screen[46][20] = 16'b11010_100100_00110;
end_screen[46][21] = 16'b11011_101110_01111;
end_screen[46][22] = 16'b11100_110010_10010;
end_screen[46][23] = 16'b11101_110101_10100;
end_screen[46][24] = 16'b11101_110100_10011;
end_screen[46][25] = 16'b11100_110011_10010;
end_screen[46][26] = 16'b11101_110101_10100;
end_screen[46][27] = 16'b11110_110110_10100;
end_screen[46][28] = 16'b11100_110010_10010;
end_screen[46][29] = 16'b11100_110010_10010;
end_screen[46][30] = 16'b11101_110101_10011;
end_screen[46][31] = 16'b11101_110100_10011;
end_screen[46][32] = 16'b11010_101010_01101;
end_screen[46][33] = 16'b11001_101000_01011;
end_screen[46][34] = 16'b11100_110001_10001;
end_screen[46][35] = 16'b11100_110001_10010;
end_screen[46][36] = 16'b10001_101010_11100;
end_screen[46][37] = 16'b10001_101010_11100;
end_screen[46][38] = 16'b10001_101010_11100;
end_screen[46][39] = 16'b11111_110011_00111;
end_screen[46][40] = 16'b11111_110011_00111;
end_screen[46][41] = 16'b11111_110011_00111;
end_screen[46][42] = 16'b11111_110011_00111;
end_screen[46][43] = 16'b11111_110011_00111;
end_screen[46][44] = 16'b11111_110011_00111;
end_screen[46][45] = 16'b11111_110011_00111;
end_screen[46][46] = 16'b11111_110011_00111;
end_screen[46][47] = 16'b11111_110011_00111;
end_screen[46][48] = 16'b11111_110011_00111;
end_screen[46][49] = 16'b11111_110011_00111;
end_screen[46][50] = 16'b11111_110011_00111;
end_screen[46][51] = 16'b11111_110011_00111;
end_screen[46][52] = 16'b11111_110011_00111;
end_screen[46][53] = 16'b11111_110011_00111;
end_screen[46][54] = 16'b11111_110011_00111;
end_screen[46][55] = 16'b11111_110011_00111;
end_screen[46][56] = 16'b11111_110011_00111;
end_screen[46][57] = 16'b11111_110011_00111;
end_screen[46][58] = 16'b10001_101010_11100;
end_screen[46][59] = 16'b10001_101010_11100;
end_screen[46][60] = 16'b10001_101010_11100;
end_screen[46][61] = 16'b10001_101010_11100;
end_screen[46][62] = 16'b10001_101010_11100;
end_screen[46][63] = 16'b10100_101011_11001;
end_screen[46][64] = 16'b11000_101100_10011;
end_screen[46][65] = 16'b11010_101110_01111;
end_screen[46][66] = 16'b11010_101000_01100;
end_screen[46][67] = 16'b10111_010000_00010;
end_screen[46][68] = 16'b10110_000101_00000;
end_screen[46][69] = 16'b10110_000111_00000;
end_screen[46][70] = 16'b11000_001101_00001;
end_screen[46][71] = 16'b11000_001110_00001;
end_screen[46][72] = 16'b11000_001101_00001;
end_screen[46][73] = 16'b11001_001111_00001;
end_screen[46][74] = 16'b11001_001111_00010;
end_screen[46][75] = 16'b11001_001110_00001;
end_screen[46][76] = 16'b11000_001110_00001;
end_screen[46][77] = 16'b11001_001111_00001;
end_screen[46][78] = 16'b11000_001110_00001;
end_screen[46][79] = 16'b11000_001101_00001;
end_screen[46][80] = 16'b11000_001101_00001;
end_screen[46][81] = 16'b11000_001101_00001;
end_screen[46][82] = 16'b11000_001101_00001;
end_screen[46][83] = 16'b11000_001100_00001;
end_screen[46][84] = 16'b11000_001100_00001;
end_screen[46][85] = 16'b10111_001100_00001;
end_screen[46][86] = 16'b11000_001110_00001;
end_screen[46][87] = 16'b11001_001111_00010;
end_screen[46][88] = 16'b11000_001010_00000;
end_screen[46][89] = 16'b10111_001000_00000;
end_screen[46][90] = 16'b11000_010100_00011;
end_screen[46][91] = 16'b11010_100110_01100;
end_screen[46][92] = 16'b11011_110001_10011;
end_screen[46][93] = 16'b11010_101100_01110;
end_screen[46][94] = 16'b10110_101000_10010;
end_screen[46][95] = 16'b10001_101010_11100;
end_screen[47][0] = 16'b10001_101010_11100;
end_screen[47][1] = 16'b11001_110000_10101;
end_screen[47][2] = 16'b11101_110011_10010;
end_screen[47][3] = 16'b11100_110011_10010;
end_screen[47][4] = 16'b11001_100110_01011;
end_screen[47][5] = 16'b10101_010100_00000;
end_screen[47][6] = 16'b10110_010111_00001;
end_screen[47][7] = 16'b10110_010101_00000;
end_screen[47][8] = 16'b11000_011010_00001;
end_screen[47][9] = 16'b11100_100100_00011;
end_screen[47][10] = 16'b11110_101001_00110;
end_screen[47][11] = 16'b11110_101011_00111;
end_screen[47][12] = 16'b11100_100111_00101;
end_screen[47][13] = 16'b11010_011110_00001;
end_screen[47][14] = 16'b11001_011101_00001;
end_screen[47][15] = 16'b11001_011110_00011;
end_screen[47][16] = 16'b11011_100101_00110;
end_screen[47][17] = 16'b11100_100111_00110;
end_screen[47][18] = 16'b11011_100101_00110;
end_screen[47][19] = 16'b11011_100100_00101;
end_screen[47][20] = 16'b11010_100010_00101;
end_screen[47][21] = 16'b11010_101011_01101;
end_screen[47][22] = 16'b11100_110001_10001;
end_screen[47][23] = 16'b11101_110011_10010;
end_screen[47][24] = 16'b11100_110010_10010;
end_screen[47][25] = 16'b11101_110011_10010;
end_screen[47][26] = 16'b11101_110100_10011;
end_screen[47][27] = 16'b11101_110011_10010;
end_screen[47][28] = 16'b11101_110101_10100;
end_screen[47][29] = 16'b11101_110101_10011;
end_screen[47][30] = 16'b11101_110100_10011;
end_screen[47][31] = 16'b11100_110010_10001;
end_screen[47][32] = 16'b11001_101000_01100;
end_screen[47][33] = 16'b11001_101000_01100;
end_screen[47][34] = 16'b11100_110010_10001;
end_screen[47][35] = 16'b11100_110001_10010;
end_screen[47][36] = 16'b10001_101010_11100;
end_screen[47][37] = 16'b10001_101010_11100;
end_screen[47][38] = 16'b10001_101010_11100;
end_screen[47][39] = 16'b11111_110011_00111;
end_screen[47][40] = 16'b11111_110011_00111;
end_screen[47][41] = 16'b11111_110011_00111;
end_screen[47][42] = 16'b11111_110011_00111;
end_screen[47][43] = 16'b11111_110011_00111;
end_screen[47][44] = 16'b11111_110011_00111;
end_screen[47][45] = 16'b11111_110011_00111;
end_screen[47][46] = 16'b11111_110011_00111;
end_screen[47][47] = 16'b11111_110011_00111;
end_screen[47][48] = 16'b11111_110011_00111;
end_screen[47][49] = 16'b11111_110011_00111;
end_screen[47][50] = 16'b11111_110011_00111;
end_screen[47][51] = 16'b11111_110011_00111;
end_screen[47][52] = 16'b11111_110011_00111;
end_screen[47][53] = 16'b11111_110011_00111;
end_screen[47][54] = 16'b11111_110011_00111;
end_screen[47][55] = 16'b11111_110011_00111;
end_screen[47][56] = 16'b11111_110011_00111;
end_screen[47][57] = 16'b11111_110011_00111;
end_screen[47][58] = 16'b10001_101010_11100;
end_screen[47][59] = 16'b10001_101010_11100;
end_screen[47][60] = 16'b10001_101010_11100;
end_screen[47][61] = 16'b10001_101010_11100;
end_screen[47][62] = 16'b10001_101010_11100;
end_screen[47][63] = 16'b10001_101010_11100;
end_screen[47][64] = 16'b10101_101010_10110;
end_screen[47][65] = 16'b11001_101001_01101;
end_screen[47][66] = 16'b11010_101111_10000;
end_screen[47][67] = 16'b11010_101000_01101;
end_screen[47][68] = 16'b11000_011000_00110;
end_screen[47][69] = 16'b10111_001101_00001;
end_screen[47][70] = 16'b10110_000110_00000;
end_screen[47][71] = 16'b10110_000110_00000;
end_screen[47][72] = 16'b10111_001010_00000;
end_screen[47][73] = 16'b11000_001101_00001;
end_screen[47][74] = 16'b11000_001101_00001;
end_screen[47][75] = 16'b11000_001101_00001;
end_screen[47][76] = 16'b11000_001101_00001;
end_screen[47][77] = 16'b11000_001110_00001;
end_screen[47][78] = 16'b11001_001111_00010;
end_screen[47][79] = 16'b11001_001111_00010;
end_screen[47][80] = 16'b11001_001110_00001;
end_screen[47][81] = 16'b11001_001110_00001;
end_screen[47][82] = 16'b11001_010000_00010;
end_screen[47][83] = 16'b11001_001111_00001;
end_screen[47][84] = 16'b11000_001110_00001;
end_screen[47][85] = 16'b11001_001110_00001;
end_screen[47][86] = 16'b11000_001010_00000;
end_screen[47][87] = 16'b10111_001000_00000;
end_screen[47][88] = 16'b10111_001101_00001;
end_screen[47][89] = 16'b11000_011001_00110;
end_screen[47][90] = 16'b11010_101100_01111;
end_screen[47][91] = 16'b11100_110100_10100;
end_screen[47][92] = 16'b11010_101011_01111;
end_screen[47][93] = 16'b10111_101000_01111;
end_screen[47][94] = 16'b10100_101010_10111;
end_screen[47][95] = 16'b10001_101010_11100;
end_screen[48][0] = 16'b10001_101010_11100;
end_screen[48][1] = 16'b11001_110001_10101;
end_screen[48][2] = 16'b11100_110010_10010;
end_screen[48][3] = 16'b11100_110010_10010;
end_screen[48][4] = 16'b11011_101101_01111;
end_screen[48][5] = 16'b10111_011111_00111;
end_screen[48][6] = 16'b10101_010110_00001;
end_screen[48][7] = 16'b11001_011100_00001;
end_screen[48][8] = 16'b11100_100100_00100;
end_screen[48][9] = 16'b11101_100111_00101;
end_screen[48][10] = 16'b11011_100000_00010;
end_screen[48][11] = 16'b10111_011000_00000;
end_screen[48][12] = 16'b11000_011001_00000;
end_screen[48][13] = 16'b11010_011101_00000;
end_screen[48][14] = 16'b11010_011111_00001;
end_screen[48][15] = 16'b11100_100111_00111;
end_screen[48][16] = 16'b11100_101001_01000;
end_screen[48][17] = 16'b11100_100101_00101;
end_screen[48][18] = 16'b11011_100100_00100;
end_screen[48][19] = 16'b11010_011111_00001;
end_screen[48][20] = 16'b11001_011110_00010;
end_screen[48][21] = 16'b11011_101110_01111;
end_screen[48][22] = 16'b11101_110100_10011;
end_screen[48][23] = 16'b11100_110001_10001;
end_screen[48][24] = 16'b11011_101110_01111;
end_screen[48][25] = 16'b11100_110001_10001;
end_screen[48][26] = 16'b11101_110100_10011;
end_screen[48][27] = 16'b11100_110010_10010;
end_screen[48][28] = 16'b11100_110010_10010;
end_screen[48][29] = 16'b11101_110011_10010;
end_screen[48][30] = 16'b11101_110100_10010;
end_screen[48][31] = 16'b11010_101100_01110;
end_screen[48][32] = 16'b11001_100111_01011;
end_screen[48][33] = 16'b11011_101101_01110;
end_screen[48][34] = 16'b11100_110010_10001;
end_screen[48][35] = 16'b11100_110001_10010;
end_screen[48][36] = 16'b10001_101010_11100;
end_screen[48][37] = 16'b10001_101010_11100;
end_screen[48][38] = 16'b10001_101010_11100;
end_screen[48][39] = 16'b11111_110011_00111;
end_screen[48][40] = 16'b11111_110011_00111;
end_screen[48][41] = 16'b11111_110011_00111;
end_screen[48][42] = 16'b11111_110011_00111;
end_screen[48][43] = 16'b11111_110011_00111;
end_screen[48][44] = 16'b11111_110011_00111;
end_screen[48][45] = 16'b11111_110011_00111;
end_screen[48][46] = 16'b11111_110011_00111;
end_screen[48][47] = 16'b11111_110011_00111;
end_screen[48][48] = 16'b11111_110011_00111;
end_screen[48][49] = 16'b11111_110011_00111;
end_screen[48][50] = 16'b11111_110011_00111;
end_screen[48][51] = 16'b11111_110011_00111;
end_screen[48][52] = 16'b11111_110011_00111;
end_screen[48][53] = 16'b11111_110011_00111;
end_screen[48][54] = 16'b11111_110011_00111;
end_screen[48][55] = 16'b11111_110011_00111;
end_screen[48][56] = 16'b11111_110011_00111;
end_screen[48][57] = 16'b11111_110011_00111;
end_screen[48][58] = 16'b10001_101010_11100;
end_screen[48][59] = 16'b10001_101010_11100;
end_screen[48][60] = 16'b10001_101010_11100;
end_screen[48][61] = 16'b10001_101010_11100;
end_screen[48][62] = 16'b10001_101010_11100;
end_screen[48][63] = 16'b10001_101010_11100;
end_screen[48][64] = 16'b10100_101010_10111;
end_screen[48][65] = 16'b11000_101000_01110;
end_screen[48][66] = 16'b11010_101010_01110;
end_screen[48][67] = 16'b11011_110001_10010;
end_screen[48][68] = 16'b11011_110011_10010;
end_screen[48][69] = 16'b11001_100011_01010;
end_screen[48][70] = 16'b11000_010100_00100;
end_screen[48][71] = 16'b10111_001110_00010;
end_screen[48][72] = 16'b10110_001011_00000;
end_screen[48][73] = 16'b10110_001000_00000;
end_screen[48][74] = 16'b10110_001000_00000;
end_screen[48][75] = 16'b10111_001001_00000;
end_screen[48][76] = 16'b10111_001011_00000;
end_screen[48][77] = 16'b11000_001100_00001;
end_screen[48][78] = 16'b11000_001101_00001;
end_screen[48][79] = 16'b11001_001101_00001;
end_screen[48][80] = 16'b11000_001100_00001;
end_screen[48][81] = 16'b11000_001011_00000;
end_screen[48][82] = 16'b11000_001011_00000;
end_screen[48][83] = 16'b10111_001010_00000;
end_screen[48][84] = 16'b10111_001001_00000;
end_screen[48][85] = 16'b11000_001011_00000;
end_screen[48][86] = 16'b11000_001111_00010;
end_screen[48][87] = 16'b11000_010110_00101;
end_screen[48][88] = 16'b11001_100100_01011;
end_screen[48][89] = 16'b11011_110010_10010;
end_screen[48][90] = 16'b11011_110010_10011;
end_screen[48][91] = 16'b11001_101010_01110;
end_screen[48][92] = 16'b11000_100111_01011;
end_screen[48][93] = 16'b10101_101011_10111;
end_screen[48][94] = 16'b10001_101010_11100;
end_screen[48][95] = 16'b10001_101010_11100;
end_screen[49][0] = 16'b10001_101010_11100;
end_screen[49][1] = 16'b11010_101111_10010;
end_screen[49][2] = 16'b11100_110001_10001;
end_screen[49][3] = 16'b11100_110010_10010;
end_screen[49][4] = 16'b11011_110000_10000;
end_screen[49][5] = 16'b11001_100111_01010;
end_screen[49][6] = 16'b10111_011011_00010;
end_screen[49][7] = 16'b11011_100000_00010;
end_screen[49][8] = 16'b11100_100010_00010;
end_screen[49][9] = 16'b11001_011101_00001;
end_screen[49][10] = 16'b10110_010100_00000;
end_screen[49][11] = 16'b10110_010110_00000;
end_screen[49][12] = 16'b11011_100010_00100;
end_screen[49][13] = 16'b11100_101000_00111;
end_screen[49][14] = 16'b11101_101011_01001;
end_screen[49][15] = 16'b11101_101101_01011;
end_screen[49][16] = 16'b11100_101010_01000;
end_screen[49][17] = 16'b11011_100011_00101;
end_screen[49][18] = 16'b11010_100000_00011;
end_screen[49][19] = 16'b11000_011011_00000;
end_screen[49][20] = 16'b10111_011110_00101;
end_screen[49][21] = 16'b11011_101101_01110;
end_screen[49][22] = 16'b11100_110010_10001;
end_screen[49][23] = 16'b11101_110011_10010;
end_screen[49][24] = 16'b11100_101111_10000;
end_screen[49][25] = 16'b11011_101111_01111;
end_screen[49][26] = 16'b11100_110001_10001;
end_screen[49][27] = 16'b11101_110011_10010;
end_screen[49][28] = 16'b11100_110010_10001;
end_screen[49][29] = 16'b11100_110010_10001;
end_screen[49][30] = 16'b11100_110000_10000;
end_screen[49][31] = 16'b11000_100100_01001;
end_screen[49][32] = 16'b11000_100101_01010;
end_screen[49][33] = 16'b11100_110001_10001;
end_screen[49][34] = 16'b11100_110010_10001;
end_screen[49][35] = 16'b11100_110001_10001;
end_screen[49][36] = 16'b10001_101010_11100;
end_screen[49][37] = 16'b10001_101010_11100;
end_screen[49][38] = 16'b10001_101010_11100;
end_screen[49][39] = 16'b11111_110011_00111;
end_screen[49][40] = 16'b11111_110011_00111;
end_screen[49][41] = 16'b11111_110011_00111;
end_screen[49][42] = 16'b11111_110011_00111;
end_screen[49][43] = 16'b11111_110011_00111;
end_screen[49][44] = 16'b11111_110011_00111;
end_screen[49][45] = 16'b11111_110011_00111;
end_screen[49][46] = 16'b11111_110011_00111;
end_screen[49][47] = 16'b11111_110011_00111;
end_screen[49][48] = 16'b11111_110011_00111;
end_screen[49][49] = 16'b11111_110011_00111;
end_screen[49][50] = 16'b11111_110011_00111;
end_screen[49][51] = 16'b11111_110011_00111;
end_screen[49][52] = 16'b11111_110011_00111;
end_screen[49][53] = 16'b11111_110011_00111;
end_screen[49][54] = 16'b11111_110011_00111;
end_screen[49][55] = 16'b11111_110011_00111;
end_screen[49][56] = 16'b11111_110011_00111;
end_screen[49][57] = 16'b11111_110011_00111;
end_screen[49][58] = 16'b10001_101010_11100;
end_screen[49][59] = 16'b10001_101010_11100;
end_screen[49][60] = 16'b10001_101010_11100;
end_screen[49][61] = 16'b10001_101010_11100;
end_screen[49][62] = 16'b10001_101010_11100;
end_screen[49][63] = 16'b10001_101010_11100;
end_screen[49][64] = 16'b10001_101010_11100;
end_screen[49][65] = 16'b10100_101011_11000;
end_screen[49][66] = 16'b11001_101000_01100;
end_screen[49][67] = 16'b11001_101001_01101;
end_screen[49][68] = 16'b11010_101100_01111;
end_screen[49][69] = 16'b11011_101111_10000;
end_screen[49][70] = 16'b11011_110010_10010;
end_screen[49][71] = 16'b11010_101100_01110;
end_screen[49][72] = 16'b11000_011100_00111;
end_screen[49][73] = 16'b10111_010001_00011;
end_screen[49][74] = 16'b10111_001110_00010;
end_screen[49][75] = 16'b10111_001101_00010;
end_screen[49][76] = 16'b10111_001100_00001;
end_screen[49][77] = 16'b10111_001011_00000;
end_screen[49][78] = 16'b10111_001011_00000;
end_screen[49][79] = 16'b10111_001011_00000;
end_screen[49][80] = 16'b10111_001010_00000;
end_screen[49][81] = 16'b10111_001011_00000;
end_screen[49][82] = 16'b10111_001100_00001;
end_screen[49][83] = 16'b10111_001101_00010;
end_screen[49][84] = 16'b10111_001011_00001;
end_screen[49][85] = 16'b11000_010100_00011;
end_screen[49][86] = 16'b11010_101001_01101;
end_screen[49][87] = 16'b11100_110100_10100;
end_screen[49][88] = 16'b11011_110010_10011;
end_screen[49][89] = 16'b11011_101110_10001;
end_screen[49][90] = 16'b11001_101001_01101;
end_screen[49][91] = 16'b11001_101001_01101;
end_screen[49][92] = 16'b11000_101001_01110;
end_screen[49][93] = 16'b10100_101010_10111;
end_screen[49][94] = 16'b10001_101010_11100;
end_screen[49][95] = 16'b10001_101010_11100;
end_screen[50][0] = 16'b10001_101010_11100;
end_screen[50][1] = 16'b10101_101100_11000;
end_screen[50][2] = 16'b11001_110000_10100;
end_screen[50][3] = 16'b11100_110010_10001;
end_screen[50][4] = 16'b11100_110001_10001;
end_screen[50][5] = 16'b11010_101011_01101;
end_screen[50][6] = 16'b11000_100001_00111;
end_screen[50][7] = 16'b11000_011011_00001;
end_screen[50][8] = 16'b11000_011001_00000;
end_screen[50][9] = 16'b11000_011000_00000;
end_screen[50][10] = 16'b11001_011011_00001;
end_screen[50][11] = 16'b11100_100100_00011;
end_screen[50][12] = 16'b11101_101010_00110;
end_screen[50][13] = 16'b11101_101010_01000;
end_screen[50][14] = 16'b11110_101101_01010;
end_screen[50][15] = 16'b11101_101100_01010;
end_screen[50][16] = 16'b11011_100101_00111;
end_screen[50][17] = 16'b11010_100100_00111;
end_screen[50][18] = 16'b11011_101000_01000;
end_screen[50][19] = 16'b11010_100100_00111;
end_screen[50][20] = 16'b10111_100010_01001;
end_screen[50][21] = 16'b11011_101100_01110;
end_screen[50][22] = 16'b11100_110000_10000;
end_screen[50][23] = 16'b11101_110011_10010;
end_screen[50][24] = 16'b11100_110010_10001;
end_screen[50][25] = 16'b11100_101111_10000;
end_screen[50][26] = 16'b11100_110001_10001;
end_screen[50][27] = 16'b11101_110011_10010;
end_screen[50][28] = 16'b11100_110010_10001;
end_screen[50][29] = 16'b11100_110001_10001;
end_screen[50][30] = 16'b11001_100111_01011;
end_screen[50][31] = 16'b10111_100010_01000;
end_screen[50][32] = 16'b11010_101010_01101;
end_screen[50][33] = 16'b11100_110001_10001;
end_screen[50][34] = 16'b11011_110000_10011;
end_screen[50][35] = 16'b10110_101101_10111;
end_screen[50][36] = 16'b10001_101010_11100;
end_screen[50][37] = 16'b10001_101010_11100;
end_screen[50][38] = 16'b10001_101010_11100;
end_screen[50][39] = 16'b11111_111111_11111;
end_screen[50][40] = 16'b11111_111111_11111;
end_screen[50][41] = 16'b11111_111111_11111;
end_screen[50][42] = 16'b11111_111111_11111;
end_screen[50][43] = 16'b11111_111111_11111;
end_screen[50][44] = 16'b11111_111111_11111;
end_screen[50][45] = 16'b01111_011110_01111;
end_screen[50][46] = 16'b01111_011110_01111;
end_screen[50][47] = 16'b01111_011110_01111;
end_screen[50][48] = 16'b01111_011110_01111;
end_screen[50][49] = 16'b01111_011110_01111;
end_screen[50][50] = 16'b01111_011110_01111;
end_screen[50][51] = 16'b01111_011110_01111;
end_screen[50][52] = 16'b11111_111111_11111;
end_screen[50][53] = 16'b11111_111111_11111;
end_screen[50][54] = 16'b11111_111111_11111;
end_screen[50][55] = 16'b11111_111111_11111;
end_screen[50][56] = 16'b11111_111111_11111;
end_screen[50][57] = 16'b11111_111111_11111;
end_screen[50][58] = 16'b10001_101010_11100;
end_screen[50][59] = 16'b10001_101010_11100;
end_screen[50][60] = 16'b10001_101010_11100;
end_screen[50][61] = 16'b10001_101010_11100;
end_screen[50][62] = 16'b10001_101010_11100;
end_screen[50][63] = 16'b10001_101010_11100;
end_screen[50][64] = 16'b10001_101010_11100;
end_screen[50][65] = 16'b10100_101011_11001;
end_screen[50][66] = 16'b11000_101000_01101;
end_screen[50][67] = 16'b11001_101001_01101;
end_screen[50][68] = 16'b11001_101000_01101;
end_screen[50][69] = 16'b11001_101001_01101;
end_screen[50][70] = 16'b11010_101101_01111;
end_screen[50][71] = 16'b11011_110000_10001;
end_screen[50][72] = 16'b11011_101111_10001;
end_screen[50][73] = 16'b11010_101100_01111;
end_screen[50][74] = 16'b11010_101011_01110;
end_screen[50][75] = 16'b11010_101001_01110;
end_screen[50][76] = 16'b11001_100000_01000;
end_screen[50][77] = 16'b11000_011001_00101;
end_screen[50][78] = 16'b10111_010111_00101;
end_screen[50][79] = 16'b10111_010111_00101;
end_screen[50][80] = 16'b11000_011001_00110;
end_screen[50][81] = 16'b11000_011101_00111;
end_screen[50][82] = 16'b11001_100100_01010;
end_screen[50][83] = 16'b11010_101011_01111;
end_screen[50][84] = 16'b11010_101011_01111;
end_screen[50][85] = 16'b11010_101011_01111;
end_screen[50][86] = 16'b11011_101110_10000;
end_screen[50][87] = 16'b11010_101101_01111;
end_screen[50][88] = 16'b11001_101001_01101;
end_screen[50][89] = 16'b11001_101001_01101;
end_screen[50][90] = 16'b11001_101001_01101;
end_screen[50][91] = 16'b11001_101001_01101;
end_screen[50][92] = 16'b10100_101011_11000;
end_screen[50][93] = 16'b10001_101010_11100;
end_screen[50][94] = 16'b10001_101010_11100;
end_screen[50][95] = 16'b10001_101010_11100;
end_screen[51][0] = 16'b10001_101010_11100;
end_screen[51][1] = 16'b10001_101010_11100;
end_screen[51][2] = 16'b10111_101111_10111;
end_screen[51][3] = 16'b11100_110001_10000;
end_screen[51][4] = 16'b11100_110011_10010;
end_screen[51][5] = 16'b11100_110001_10001;
end_screen[51][6] = 16'b11001_100111_01011;
end_screen[51][7] = 16'b10110_011100_00100;
end_screen[51][8] = 16'b10101_010111_00010;
end_screen[51][9] = 16'b11001_011011_00001;
end_screen[51][10] = 16'b11101_100100_00010;
end_screen[51][11] = 16'b11101_100110_00100;
end_screen[51][12] = 16'b11011_100010_00011;
end_screen[51][13] = 16'b11100_100011_00011;
end_screen[51][14] = 16'b11011_100010_00011;
end_screen[51][15] = 16'b11011_100101_00110;
end_screen[51][16] = 16'b11010_100101_01000;
end_screen[51][17] = 16'b11011_101001_01011;
end_screen[51][18] = 16'b11100_101011_01011;
end_screen[51][19] = 16'b11001_100011_00111;
end_screen[51][20] = 16'b11000_100100_01001;
end_screen[51][21] = 16'b11011_101101_01110;
end_screen[51][22] = 16'b11101_110010_10001;
end_screen[51][23] = 16'b11100_110000_10000;
end_screen[51][24] = 16'b11011_101101_01111;
end_screen[51][25] = 16'b11100_110000_10000;
end_screen[51][26] = 16'b11101_110011_10010;
end_screen[51][27] = 16'b11100_110000_10000;
end_screen[51][28] = 16'b11010_101001_01100;
end_screen[51][29] = 16'b11001_100111_01011;
end_screen[51][30] = 16'b10111_100010_01000;
end_screen[51][31] = 16'b11010_101001_01100;
end_screen[51][32] = 16'b11100_110001_10001;
end_screen[51][33] = 16'b11100_101111_10000;
end_screen[51][34] = 16'b11001_101110_10010;
end_screen[51][35] = 16'b10001_101010_11100;
end_screen[51][36] = 16'b10001_101010_11100;
end_screen[51][37] = 16'b10001_101010_11100;
end_screen[51][38] = 16'b10001_101010_11100;
end_screen[51][39] = 16'b11111_111111_11111;
end_screen[51][40] = 16'b11111_111111_11111;
end_screen[51][41] = 16'b11111_111111_11111;
end_screen[51][42] = 16'b11111_111111_11111;
end_screen[51][43] = 16'b11111_111111_11111;
end_screen[51][44] = 16'b11111_111111_11111;
end_screen[51][45] = 16'b01111_011110_01111;
end_screen[51][46] = 16'b01111_011110_01111;
end_screen[51][47] = 16'b01110_011101_01111;
end_screen[51][48] = 16'b01110_011101_01111;
end_screen[51][49] = 16'b01110_011101_01111;
end_screen[51][50] = 16'b01111_011110_01111;
end_screen[51][51] = 16'b01111_011110_01111;
end_screen[51][52] = 16'b11111_111111_11111;
end_screen[51][53] = 16'b11111_111111_11111;
end_screen[51][54] = 16'b11111_111111_11111;
end_screen[51][55] = 16'b11111_111111_11111;
end_screen[51][56] = 16'b11111_111111_11111;
end_screen[51][57] = 16'b11111_111111_11111;
end_screen[51][58] = 16'b10001_101010_11100;
end_screen[51][59] = 16'b10001_101010_11100;
end_screen[51][60] = 16'b10001_101010_11100;
end_screen[51][61] = 16'b10001_101010_11100;
end_screen[51][62] = 16'b10001_101010_11100;
end_screen[51][63] = 16'b10001_101010_11100;
end_screen[51][64] = 16'b10001_101010_11100;
end_screen[51][65] = 16'b10001_101010_11100;
end_screen[51][66] = 16'b10011_101010_11001;
end_screen[51][67] = 16'b11001_101010_01101;
end_screen[51][68] = 16'b11001_101001_01101;
end_screen[51][69] = 16'b11001_101001_01101;
end_screen[51][70] = 16'b11001_101001_01101;
end_screen[51][71] = 16'b11001_101010_01110;
end_screen[51][72] = 16'b11010_101100_01111;
end_screen[51][73] = 16'b11010_101101_01111;
end_screen[51][74] = 16'b11010_101110_01111;
end_screen[51][75] = 16'b11011_110000_10001;
end_screen[51][76] = 16'b11011_110000_10001;
end_screen[51][77] = 16'b11010_101101_10000;
end_screen[51][78] = 16'b11010_101011_01110;
end_screen[51][79] = 16'b11010_101011_01110;
end_screen[51][80] = 16'b11010_101100_01111;
end_screen[51][81] = 16'b11011_101110_10000;
end_screen[51][82] = 16'b11011_101111_10001;
end_screen[51][83] = 16'b11011_110000_10001;
end_screen[51][84] = 16'b11010_101101_01111;
end_screen[51][85] = 16'b11001_101011_01110;
end_screen[51][86] = 16'b11001_101010_01110;
end_screen[51][87] = 16'b11001_101001_01101;
end_screen[51][88] = 16'b11001_101001_01101;
end_screen[51][89] = 16'b11001_101001_01101;
end_screen[51][90] = 16'b11001_101010_01101;
end_screen[51][91] = 16'b11001_101001_01101;
end_screen[51][92] = 16'b10011_101010_11001;
end_screen[51][93] = 16'b10001_101010_11100;
end_screen[51][94] = 16'b10001_101010_11100;
end_screen[51][95] = 16'b10001_101010_11100;
end_screen[52][0] = 16'b10001_101010_11100;
end_screen[52][1] = 16'b10001_101010_11100;
end_screen[52][2] = 16'b10100_101011_10111;
end_screen[52][3] = 16'b11001_101101_10000;
end_screen[52][4] = 16'b11100_110010_10001;
end_screen[52][5] = 16'b11100_110000_10000;
end_screen[52][6] = 16'b11011_101101_01111;
end_screen[52][7] = 16'b11001_100110_01010;
end_screen[52][8] = 16'b10110_011100_00100;
end_screen[52][9] = 16'b10111_011000_00000;
end_screen[52][10] = 16'b11001_011100_00000;
end_screen[52][11] = 16'b11010_011110_00001;
end_screen[52][12] = 16'b11010_011111_00010;
end_screen[52][13] = 16'b11010_100010_00100;
end_screen[52][14] = 16'b11010_100010_00110;
end_screen[52][15] = 16'b11010_101000_01010;
end_screen[52][16] = 16'b11100_101100_01101;
end_screen[52][17] = 16'b11100_101011_01011;
end_screen[52][18] = 16'b11001_100010_00110;
end_screen[52][19] = 16'b10111_011100_00011;
end_screen[52][20] = 16'b11000_100011_01000;
end_screen[52][21] = 16'b11001_100110_01010;
end_screen[52][22] = 16'b11100_101111_01111;
end_screen[52][23] = 16'b11011_101100_01110;
end_screen[52][24] = 16'b11001_101000_01100;
end_screen[52][25] = 16'b11010_101001_01100;
end_screen[52][26] = 16'b11010_101010_01101;
end_screen[52][27] = 16'b11001_101000_01011;
end_screen[52][28] = 16'b11000_100101_01010;
end_screen[52][29] = 16'b11000_100100_01010;
end_screen[52][30] = 16'b11010_101010_01101;
end_screen[52][31] = 16'b11100_110000_10000;
end_screen[52][32] = 16'b11100_110001_10001;
end_screen[52][33] = 16'b11010_101100_01111;
end_screen[52][34] = 16'b10101_101010_10100;
end_screen[52][35] = 16'b10001_101010_11100;
end_screen[52][36] = 16'b10001_101010_11100;
end_screen[52][37] = 16'b10001_101010_11100;
end_screen[52][38] = 16'b10001_101010_11100;
end_screen[52][39] = 16'b11111_111111_11111;
end_screen[52][40] = 16'b11111_111111_11111;
end_screen[52][41] = 16'b11111_111111_11111;
end_screen[52][42] = 16'b11111_111111_11111;
end_screen[52][43] = 16'b11111_111111_11111;
end_screen[52][44] = 16'b11111_111111_11111;
end_screen[52][45] = 16'b01111_011110_01111;
end_screen[52][46] = 16'b01111_011110_01111;
end_screen[52][47] = 16'b01111_011110_01111;
end_screen[52][48] = 16'b01111_011110_01111;
end_screen[52][49] = 16'b01111_011110_01111;
end_screen[52][50] = 16'b01111_011110_01111;
end_screen[52][51] = 16'b01111_011110_01111;
end_screen[52][52] = 16'b11111_111111_11111;
end_screen[52][53] = 16'b11111_111111_11111;
end_screen[52][54] = 16'b11111_111111_11111;
end_screen[52][55] = 16'b11111_111111_11111;
end_screen[52][56] = 16'b11111_111111_11111;
end_screen[52][57] = 16'b11111_111111_11111;
end_screen[52][58] = 16'b10001_101010_11100;
end_screen[52][59] = 16'b10001_101010_11100;
end_screen[52][60] = 16'b10001_101010_11100;
end_screen[52][61] = 16'b10001_101010_11100;
end_screen[52][62] = 16'b10001_101010_11100;
end_screen[52][63] = 16'b10001_101010_11100;
end_screen[52][64] = 16'b10001_101010_11100;
end_screen[52][65] = 16'b10001_101010_11100;
end_screen[52][66] = 16'b10010_101010_11011;
end_screen[52][67] = 16'b11001_101001_01101;
end_screen[52][68] = 16'b11001_101010_01101;
end_screen[52][69] = 16'b11001_101010_01110;
end_screen[52][70] = 16'b11001_101010_01101;
end_screen[52][71] = 16'b11001_101001_01101;
end_screen[52][72] = 16'b11001_101001_01101;
end_screen[52][73] = 16'b11001_101010_01101;
end_screen[52][74] = 16'b11001_101010_01110;
end_screen[52][75] = 16'b11001_101011_01110;
end_screen[52][76] = 16'b11010_101100_01111;
end_screen[52][77] = 16'b11010_101100_01111;
end_screen[52][78] = 16'b11010_101100_01111;
end_screen[52][79] = 16'b11010_101100_01111;
end_screen[52][80] = 16'b11010_101100_01111;
end_screen[52][81] = 16'b11010_101100_01111;
end_screen[52][82] = 16'b11010_101011_01110;
end_screen[52][83] = 16'b11001_101010_01110;
end_screen[52][84] = 16'b11001_101010_01101;
end_screen[52][85] = 16'b11001_101001_01101;
end_screen[52][86] = 16'b11001_101001_01101;
end_screen[52][87] = 16'b11001_101010_01110;
end_screen[52][88] = 16'b11010_101011_01110;
end_screen[52][89] = 16'b11001_101010_01110;
end_screen[52][90] = 16'b11001_101010_01101;
end_screen[52][91] = 16'b10100_101010_11000;
end_screen[52][92] = 16'b10001_101010_11011;
end_screen[52][93] = 16'b10001_101010_11100;
end_screen[52][94] = 16'b10001_101010_11100;
end_screen[52][95] = 16'b10001_101010_11100;
end_screen[53][0] = 16'b10001_101010_11100;
end_screen[53][1] = 16'b10001_101010_11100;
end_screen[53][2] = 16'b10001_101010_11100;
end_screen[53][3] = 16'b10011_101011_11010;
end_screen[53][4] = 16'b11011_110001_10011;
end_screen[53][5] = 16'b11100_110001_10001;
end_screen[53][6] = 16'b11100_110010_10001;
end_screen[53][7] = 16'b11011_101101_01111;
end_screen[53][8] = 16'b11000_100011_01001;
end_screen[53][9] = 16'b10110_011011_00100;
end_screen[53][10] = 16'b10101_011000_00010;
end_screen[53][11] = 16'b10111_011001_00001;
end_screen[53][12] = 16'b11001_011111_00011;
end_screen[53][13] = 16'b11011_100110_00111;
end_screen[53][14] = 16'b11101_101100_01100;
end_screen[53][15] = 16'b11101_110001_10001;
end_screen[53][16] = 16'b11100_101101_01101;
end_screen[53][17] = 16'b11001_100010_00110;
end_screen[53][18] = 16'b10111_011011_00011;
end_screen[53][19] = 16'b10110_011011_00100;
end_screen[53][20] = 16'b10111_100001_00111;
end_screen[53][21] = 16'b10111_100010_01000;
end_screen[53][22] = 16'b11001_100111_01011;
end_screen[53][23] = 16'b11001_101000_01011;
end_screen[53][24] = 16'b11001_100111_01011;
end_screen[53][25] = 16'b11000_100100_01001;
end_screen[53][26] = 16'b11000_100011_01001;
end_screen[53][27] = 16'b11001_100111_01011;
end_screen[53][28] = 16'b11010_101011_01101;
end_screen[53][29] = 16'b11100_110000_10000;
end_screen[53][30] = 16'b11100_110001_10001;
end_screen[53][31] = 16'b11100_110000_10000;
end_screen[53][32] = 16'b11011_110000_10001;
end_screen[53][33] = 16'b10110_101101_10111;
end_screen[53][34] = 16'b10001_101010_11100;
end_screen[53][35] = 16'b10001_101010_11100;
end_screen[53][36] = 16'b10001_101010_11100;
end_screen[53][37] = 16'b10001_101010_11100;
end_screen[53][38] = 16'b10001_101010_11100;
end_screen[53][39] = 16'b11111_111111_11111;
end_screen[53][40] = 16'b11111_111111_11111;
end_screen[53][41] = 16'b11111_111111_11111;
end_screen[53][42] = 16'b11111_111111_11111;
end_screen[53][43] = 16'b11111_111111_11111;
end_screen[53][44] = 16'b11111_111111_11111;
end_screen[53][45] = 16'b10010_100101_10010;
end_screen[53][46] = 16'b10010_100101_10010;
end_screen[53][47] = 16'b10010_100101_10010;
end_screen[53][48] = 16'b10010_100101_10010;
end_screen[53][49] = 16'b10010_100101_10010;
end_screen[53][50] = 16'b10010_100101_10010;
end_screen[53][51] = 16'b10010_100101_10010;
end_screen[53][52] = 16'b11111_111111_11111;
end_screen[53][53] = 16'b11111_111111_11111;
end_screen[53][54] = 16'b11111_111111_11111;
end_screen[53][55] = 16'b11111_111111_11111;
end_screen[53][56] = 16'b11111_111111_11111;
end_screen[53][57] = 16'b11111_111111_11111;
end_screen[53][58] = 16'b10001_101010_11100;
end_screen[53][59] = 16'b10001_101010_11100;
end_screen[53][60] = 16'b10001_101010_11100;
end_screen[53][61] = 16'b10001_101010_11100;
end_screen[53][62] = 16'b10001_101010_11100;
end_screen[53][63] = 16'b10001_101010_11100;
end_screen[53][64] = 16'b10001_101010_11100;
end_screen[53][65] = 16'b10001_101010_11100;
end_screen[53][66] = 16'b10001_101010_11100;
end_screen[53][67] = 16'b10011_101011_11001;
end_screen[53][68] = 16'b11001_101001_01101;
end_screen[53][69] = 16'b11001_101010_01101;
end_screen[53][70] = 16'b11001_101010_01110;
end_screen[53][71] = 16'b11001_101010_01101;
end_screen[53][72] = 16'b11001_101010_01101;
end_screen[53][73] = 16'b11001_101010_01110;
end_screen[53][74] = 16'b11001_101010_01110;
end_screen[53][75] = 16'b11001_101001_01101;
end_screen[53][76] = 16'b11001_101001_01101;
end_screen[53][77] = 16'b11001_101001_01101;
end_screen[53][78] = 16'b11001_101010_01101;
end_screen[53][79] = 16'b11001_101001_01101;
end_screen[53][80] = 16'b11001_101001_01101;
end_screen[53][81] = 16'b11001_101001_01101;
end_screen[53][82] = 16'b11001_101001_01101;
end_screen[53][83] = 16'b11001_101001_01101;
end_screen[53][84] = 16'b11010_101011_01110;
end_screen[53][85] = 16'b11001_101011_01110;
end_screen[53][86] = 16'b11001_101010_01101;
end_screen[53][87] = 16'b11010_101011_01110;
end_screen[53][88] = 16'b11010_101011_01110;
end_screen[53][89] = 16'b11001_101001_01101;
end_screen[53][90] = 16'b10011_101011_11001;
end_screen[53][91] = 16'b10001_101010_11100;
end_screen[53][92] = 16'b10001_101010_11100;
end_screen[53][93] = 16'b10001_101010_11100;
end_screen[53][94] = 16'b10001_101010_11100;
end_screen[53][95] = 16'b10001_101010_11100;
end_screen[54][0] = 16'b10001_101010_11100;
end_screen[54][1] = 16'b10001_101010_11100;
end_screen[54][2] = 16'b10001_101010_11100;
end_screen[54][3] = 16'b10001_101010_11100;
end_screen[54][4] = 16'b10011_101011_11010;
end_screen[54][5] = 16'b11011_101110_10000;
end_screen[54][6] = 16'b11100_101111_10000;
end_screen[54][7] = 16'b11100_110000_10000;
end_screen[54][8] = 16'b11100_110001_10001;
end_screen[54][9] = 16'b11011_101101_01110;
end_screen[54][10] = 16'b11000_100010_01000;
end_screen[54][11] = 16'b10101_011011_00100;
end_screen[54][12] = 16'b10110_011110_00110;
end_screen[54][13] = 16'b11001_100011_01000;
end_screen[54][14] = 16'b11001_100001_00101;
end_screen[54][15] = 16'b11001_100010_00111;
end_screen[54][16] = 16'b11001_100011_01000;
end_screen[54][17] = 16'b10111_011110_00101;
end_screen[54][18] = 16'b10110_011100_00100;
end_screen[54][19] = 16'b11000_100011_01000;
end_screen[54][20] = 16'b11001_100110_01010;
end_screen[54][21] = 16'b11000_100101_01010;
end_screen[54][22] = 16'b11001_100110_01011;
end_screen[54][23] = 16'b11010_101001_01100;
end_screen[54][24] = 16'b11010_101001_01100;
end_screen[54][25] = 16'b11010_101100_01110;
end_screen[54][26] = 16'b11100_110000_10000;
end_screen[54][27] = 16'b11100_110001_10001;
end_screen[54][28] = 16'b11100_110001_10001;
end_screen[54][29] = 16'b11100_110001_10001;
end_screen[54][30] = 16'b11100_110000_10000;
end_screen[54][31] = 16'b11100_110001_10001;
end_screen[54][32] = 16'b10110_101101_10111;
end_screen[54][33] = 16'b10001_101010_11100;
end_screen[54][34] = 16'b10001_101010_11100;
end_screen[54][35] = 16'b10001_101010_11100;
end_screen[54][36] = 16'b10001_101010_11100;
end_screen[54][37] = 16'b10001_101010_11100;
end_screen[54][38] = 16'b10001_101010_11100;
end_screen[54][39] = 16'b11111_111111_11111;
end_screen[54][40] = 16'b11111_111111_11111;
end_screen[54][41] = 16'b11111_111111_11111;
end_screen[54][42] = 16'b11111_111111_11111;
end_screen[54][43] = 16'b11111_111111_11111;
end_screen[54][44] = 16'b11111_111111_11111;
end_screen[54][45] = 16'b10010_100101_10010;
end_screen[54][46] = 16'b10010_100100_10010;
end_screen[54][47] = 16'b10010_100101_10010;
end_screen[54][48] = 16'b10010_100101_10010;
end_screen[54][49] = 16'b10010_100101_10010;
end_screen[54][50] = 16'b10010_100101_10010;
end_screen[54][51] = 16'b10010_100101_10010;
end_screen[54][52] = 16'b11111_111111_11111;
end_screen[54][53] = 16'b11111_111111_11111;
end_screen[54][54] = 16'b11111_111111_11111;
end_screen[54][55] = 16'b11111_111111_11111;
end_screen[54][56] = 16'b11111_111111_11111;
end_screen[54][57] = 16'b11111_111111_11111;
end_screen[54][58] = 16'b10001_101010_11100;
end_screen[54][59] = 16'b10001_101010_11100;
end_screen[54][60] = 16'b10001_101010_11100;
end_screen[54][61] = 16'b10001_101010_11100;
end_screen[54][62] = 16'b10001_101010_11100;
end_screen[54][63] = 16'b10001_101010_11100;
end_screen[54][64] = 16'b10001_101010_11100;
end_screen[54][65] = 16'b10001_101010_11100;
end_screen[54][66] = 16'b10001_101010_11100;
end_screen[54][67] = 16'b10001_101010_11100;
end_screen[54][68] = 16'b10100_101011_11000;
end_screen[54][69] = 16'b11001_101010_01110;
end_screen[54][70] = 16'b11001_101001_01101;
end_screen[54][71] = 16'b11001_101010_01101;
end_screen[54][72] = 16'b11001_101011_01110;
end_screen[54][73] = 16'b11010_101011_01110;
end_screen[54][74] = 16'b11010_101011_01110;
end_screen[54][75] = 16'b11001_101011_01110;
end_screen[54][76] = 16'b11010_101011_01110;
end_screen[54][77] = 16'b11001_101011_01110;
end_screen[54][78] = 16'b11001_101010_01110;
end_screen[54][79] = 16'b11001_101010_01101;
end_screen[54][80] = 16'b11001_101010_01101;
end_screen[54][81] = 16'b11001_101010_01101;
end_screen[54][82] = 16'b11001_101010_01101;
end_screen[54][83] = 16'b11001_101010_01110;
end_screen[54][84] = 16'b11010_101100_01111;
end_screen[54][85] = 16'b11010_101011_01110;
end_screen[54][86] = 16'b11001_101010_01101;
end_screen[54][87] = 16'b11001_101001_01101;
end_screen[54][88] = 16'b11010_101010_01110;
end_screen[54][89] = 16'b10100_101010_11000;
end_screen[54][90] = 16'b10001_101010_11100;
end_screen[54][91] = 16'b10001_101010_11100;
end_screen[54][92] = 16'b10001_101010_11100;
end_screen[54][93] = 16'b10001_101010_11100;
end_screen[54][94] = 16'b10001_101010_11100;
end_screen[54][95] = 16'b10001_101010_11100;
end_screen[55][0] = 16'b10001_101010_11100;
end_screen[55][1] = 16'b10001_101010_11100;
end_screen[55][2] = 16'b10001_101010_11100;
end_screen[55][3] = 16'b10001_101010_11100;
end_screen[55][4] = 16'b10001_101010_11100;
end_screen[55][5] = 16'b10011_101010_11001;
end_screen[55][6] = 16'b11001_101000_01100;
end_screen[55][7] = 16'b11011_101110_01111;
end_screen[55][8] = 16'b11100_110001_10001;
end_screen[55][9] = 16'b11100_110000_10000;
end_screen[55][10] = 16'b11011_101101_01111;
end_screen[55][11] = 16'b11001_101001_01100;
end_screen[55][12] = 16'b11000_100110_01011;
end_screen[55][13] = 16'b11000_100011_01001;
end_screen[55][14] = 16'b10110_011111_00111;
end_screen[55][15] = 16'b10110_011110_00110;
end_screen[55][16] = 16'b10111_100000_00111;
end_screen[55][17] = 16'b11000_100010_01000;
end_screen[55][18] = 16'b11001_100111_01011;
end_screen[55][19] = 16'b11010_101100_01110;
end_screen[55][20] = 16'b11010_101011_01101;
end_screen[55][21] = 16'b11010_101100_01110;
end_screen[55][22] = 16'b11011_101110_01111;
end_screen[55][23] = 16'b11100_101111_10000;
end_screen[55][24] = 16'b11100_101111_10000;
end_screen[55][25] = 16'b11100_110001_10001;
end_screen[55][26] = 16'b11100_110001_10001;
end_screen[55][27] = 16'b11100_110001_10001;
end_screen[55][28] = 16'b11100_110001_10001;
end_screen[55][29] = 16'b11100_110001_10001;
end_screen[55][30] = 16'b11010_101011_01101;
end_screen[55][31] = 16'b10100_101001_10101;
end_screen[55][32] = 16'b10001_101010_11100;
end_screen[55][33] = 16'b10001_101010_11100;
end_screen[55][34] = 16'b10001_101010_11100;
end_screen[55][35] = 16'b10001_101010_11100;
end_screen[55][36] = 16'b10001_101010_11100;
end_screen[55][37] = 16'b10001_101010_11100;
end_screen[55][38] = 16'b10001_101010_11100;
end_screen[55][39] = 16'b11111_111111_11111;
end_screen[55][40] = 16'b11111_111111_11111;
end_screen[55][41] = 16'b11111_111111_11111;
end_screen[55][42] = 16'b11111_111111_11111;
end_screen[55][43] = 16'b11111_111111_11111;
end_screen[55][44] = 16'b11111_111111_11111;
end_screen[55][45] = 16'b10010_100101_10010;
end_screen[55][46] = 16'b10010_100101_10010;
end_screen[55][47] = 16'b10010_100101_10010;
end_screen[55][48] = 16'b10010_100101_10010;
end_screen[55][49] = 16'b10010_100101_10010;
end_screen[55][50] = 16'b10010_100101_10010;
end_screen[55][51] = 16'b10010_100101_10010;
end_screen[55][52] = 16'b11111_111111_11111;
end_screen[55][53] = 16'b11111_111111_11111;
end_screen[55][54] = 16'b11111_111111_11111;
end_screen[55][55] = 16'b11111_111111_11111;
end_screen[55][56] = 16'b11111_111111_11111;
end_screen[55][57] = 16'b11111_111111_11111;
end_screen[55][58] = 16'b10001_101010_11100;
end_screen[55][59] = 16'b10001_101010_11100;
end_screen[55][60] = 16'b10001_101010_11100;
end_screen[55][61] = 16'b10001_101010_11100;
end_screen[55][62] = 16'b10001_101010_11100;
end_screen[55][63] = 16'b10001_101010_11100;
end_screen[55][64] = 16'b10001_101010_11100;
end_screen[55][65] = 16'b10001_101010_11100;
end_screen[55][66] = 16'b10001_101010_11100;
end_screen[55][67] = 16'b10001_101010_11100;
end_screen[55][68] = 16'b10001_101010_11100;
end_screen[55][69] = 16'b10100_101010_10111;
end_screen[55][70] = 16'b10101_101010_10100;
end_screen[55][71] = 16'b11000_101010_10000;
end_screen[55][72] = 16'b11001_101010_01101;
end_screen[55][73] = 16'b11001_101010_01101;
end_screen[55][74] = 16'b11001_101010_01110;
end_screen[55][75] = 16'b11010_101011_01110;
end_screen[55][76] = 16'b11010_101011_01110;
end_screen[55][77] = 16'b11010_101011_01110;
end_screen[55][78] = 16'b11010_101011_01110;
end_screen[55][79] = 16'b11001_101010_01101;
end_screen[55][80] = 16'b11001_101010_01101;
end_screen[55][81] = 16'b11001_101010_01110;
end_screen[55][82] = 16'b11010_101011_01110;
end_screen[55][83] = 16'b11001_101010_01110;
end_screen[55][84] = 16'b11001_101010_01101;
end_screen[55][85] = 16'b11001_101001_01100;
end_screen[55][86] = 16'b11000_101010_10000;
end_screen[55][87] = 16'b10101_101011_10110;
end_screen[55][88] = 16'b10100_101010_11000;
end_screen[55][89] = 16'b10001_101010_11100;
end_screen[55][90] = 16'b10001_101010_11100;
end_screen[55][91] = 16'b10001_101010_11100;
end_screen[55][92] = 16'b10001_101010_11100;
end_screen[55][93] = 16'b10001_101010_11100;
end_screen[55][94] = 16'b10001_101010_11100;
end_screen[55][95] = 16'b10001_101010_11100;
end_screen[56][0] = 16'b10001_101010_11100;
end_screen[56][1] = 16'b10001_101010_11100;
end_screen[56][2] = 16'b10001_101010_11100;
end_screen[56][3] = 16'b10001_101010_11100;
end_screen[56][4] = 16'b10001_101010_11100;
end_screen[56][5] = 16'b10001_101010_11100;
end_screen[56][6] = 16'b10011_101001_11000;
end_screen[56][7] = 16'b11001_101001_01100;
end_screen[56][8] = 16'b11011_101110_01111;
end_screen[56][9] = 16'b11100_110001_10000;
end_screen[56][10] = 16'b11100_110000_10000;
end_screen[56][11] = 16'b11011_101111_10000;
end_screen[56][12] = 16'b11011_101101_01111;
end_screen[56][13] = 16'b11010_101100_01110;
end_screen[56][14] = 16'b11001_101001_01100;
end_screen[56][15] = 16'b11001_101010_01101;
end_screen[56][16] = 16'b11010_101011_01110;
end_screen[56][17] = 16'b11011_101101_01110;
end_screen[56][18] = 16'b11011_101101_01111;
end_screen[56][19] = 16'b11011_101110_01111;
end_screen[56][20] = 16'b11011_101111_10000;
end_screen[56][21] = 16'b11100_110000_10000;
end_screen[56][22] = 16'b11100_110001_10001;
end_screen[56][23] = 16'b11100_110000_10000;
end_screen[56][24] = 16'b11100_110001_10001;
end_screen[56][25] = 16'b11100_110010_10001;
end_screen[56][26] = 16'b11100_110001_10001;
end_screen[56][27] = 16'b11100_110000_10000;
end_screen[56][28] = 16'b11011_101110_01111;
end_screen[56][29] = 16'b10100_101011_11000;
end_screen[56][30] = 16'b10011_101010_11000;
end_screen[56][31] = 16'b10001_101010_11011;
end_screen[56][32] = 16'b10001_101010_11100;
end_screen[56][33] = 16'b10001_101010_11100;
end_screen[56][34] = 16'b10001_101010_11100;
end_screen[56][35] = 16'b10001_101010_11100;
end_screen[56][36] = 16'b10001_101010_11100;
end_screen[56][37] = 16'b10001_101010_11100;
end_screen[56][38] = 16'b10001_101010_11100;
end_screen[56][39] = 16'b11111_110011_00111;
end_screen[56][40] = 16'b11111_110011_00111;
end_screen[56][41] = 16'b11111_110011_00111;
end_screen[56][42] = 16'b11111_110011_00111;
end_screen[56][43] = 16'b10001_101010_11100;
end_screen[56][44] = 16'b10001_101010_11100;
end_screen[56][45] = 16'b10001_101010_11100;
end_screen[56][46] = 16'b10001_101010_11100;
end_screen[56][47] = 16'b10001_101010_11100;
end_screen[56][48] = 16'b10001_101010_11100;
end_screen[56][49] = 16'b10001_101010_11100;
end_screen[56][50] = 16'b10001_101010_11100;
end_screen[56][51] = 16'b10001_101010_11100;
end_screen[56][52] = 16'b10001_101010_11100;
end_screen[56][53] = 16'b10001_101010_11100;
end_screen[56][54] = 16'b11111_110011_00111;
end_screen[56][55] = 16'b11111_110011_00111;
end_screen[56][56] = 16'b11111_110011_00111;
end_screen[56][57] = 16'b11111_110011_00111;
end_screen[56][58] = 16'b10001_101010_11100;
end_screen[56][59] = 16'b10001_101010_11100;
end_screen[56][60] = 16'b10001_101010_11100;
end_screen[56][61] = 16'b10001_101010_11100;
end_screen[56][62] = 16'b10001_101010_11100;
end_screen[56][63] = 16'b10001_101010_11100;
end_screen[56][64] = 16'b10001_101010_11100;
end_screen[56][65] = 16'b10001_101010_11100;
end_screen[56][66] = 16'b10001_101010_11100;
end_screen[56][67] = 16'b10001_101010_11100;
end_screen[56][68] = 16'b10001_101010_11100;
end_screen[56][69] = 16'b10001_101010_11100;
end_screen[56][70] = 16'b10001_101010_11100;
end_screen[56][71] = 16'b10011_101010_11001;
end_screen[56][72] = 16'b10110_101001_10010;
end_screen[56][73] = 16'b10111_101001_10000;
end_screen[56][74] = 16'b11001_101001_01100;
end_screen[56][75] = 16'b11001_101001_01101;
end_screen[56][76] = 16'b11001_101000_01100;
end_screen[56][77] = 16'b11001_101001_01101;
end_screen[56][78] = 16'b11001_101010_01101;
end_screen[56][79] = 16'b11001_101000_01100;
end_screen[56][80] = 16'b11001_101000_01100;
end_screen[56][81] = 16'b11001_101001_01101;
end_screen[56][82] = 16'b11001_101001_01101;
end_screen[56][83] = 16'b11001_101001_01101;
end_screen[56][84] = 16'b10111_101010_10011;
end_screen[56][85] = 16'b10110_101010_10100;
end_screen[56][86] = 16'b10010_101010_11010;
end_screen[56][87] = 16'b10001_101010_11100;
end_screen[56][88] = 16'b10001_101010_11100;
end_screen[56][89] = 16'b10001_101010_11100;
end_screen[56][90] = 16'b10001_101010_11100;
end_screen[56][91] = 16'b10001_101010_11100;
end_screen[56][92] = 16'b10001_101010_11100;
end_screen[56][93] = 16'b10001_101010_11100;
end_screen[56][94] = 16'b10001_101010_11100;
end_screen[56][95] = 16'b10001_101010_11100;
end_screen[57][0] = 16'b10001_101010_11100;
end_screen[57][1] = 16'b10001_101010_11100;
end_screen[57][2] = 16'b10001_101010_11100;
end_screen[57][3] = 16'b10001_101010_11100;
end_screen[57][4] = 16'b10001_101010_11100;
end_screen[57][5] = 16'b10001_101010_11100;
end_screen[57][6] = 16'b10001_101010_11100;
end_screen[57][7] = 16'b10011_101001_11000;
end_screen[57][8] = 16'b10100_101010_10111;
end_screen[57][9] = 16'b10100_101100_11000;
end_screen[57][10] = 16'b11000_101011_10001;
end_screen[57][11] = 16'b11011_101100_01110;
end_screen[57][12] = 16'b11100_110001_10001;
end_screen[57][13] = 16'b11100_110000_10000;
end_screen[57][14] = 16'b11100_101111_01111;
end_screen[57][15] = 16'b11100_101111_10000;
end_screen[57][16] = 16'b11100_110001_10001;
end_screen[57][17] = 16'b11100_110010_10001;
end_screen[57][18] = 16'b11100_110000_10000;
end_screen[57][19] = 16'b11100_110000_10000;
end_screen[57][20] = 16'b11100_110001_10001;
end_screen[57][21] = 16'b11100_110001_10001;
end_screen[57][22] = 16'b11100_110010_10001;
end_screen[57][23] = 16'b11100_110001_10001;
end_screen[57][24] = 16'b11100_110001_10001;
end_screen[57][25] = 16'b11011_101111_10000;
end_screen[57][26] = 16'b11010_101110_10001;
end_screen[57][27] = 16'b10100_101100_11000;
end_screen[57][28] = 16'b10100_101010_10111;
end_screen[57][29] = 16'b10001_101010_11100;
end_screen[57][30] = 16'b10001_101010_11100;
end_screen[57][31] = 16'b10001_101010_11100;
end_screen[57][32] = 16'b10001_101010_11100;
end_screen[57][33] = 16'b10001_101010_11100;
end_screen[57][34] = 16'b10001_101010_11100;
end_screen[57][35] = 16'b10001_101010_11100;
end_screen[57][36] = 16'b10001_101010_11100;
end_screen[57][37] = 16'b10001_101010_11100;
end_screen[57][38] = 16'b10001_101010_11100;
end_screen[57][39] = 16'b11111_110011_00111;
end_screen[57][40] = 16'b11111_110011_00111;
end_screen[57][41] = 16'b11111_110011_00111;
end_screen[57][42] = 16'b11111_110011_00111;
end_screen[57][43] = 16'b10001_101010_11100;
end_screen[57][44] = 16'b10001_101010_11100;
end_screen[57][45] = 16'b10001_101010_11100;
end_screen[57][46] = 16'b10001_101010_11100;
end_screen[57][47] = 16'b10001_101010_11100;
end_screen[57][48] = 16'b10001_101010_11100;
end_screen[57][49] = 16'b10001_101010_11100;
end_screen[57][50] = 16'b10001_101010_11100;
end_screen[57][51] = 16'b10001_101010_11100;
end_screen[57][52] = 16'b10001_101010_11100;
end_screen[57][53] = 16'b10001_101010_11100;
end_screen[57][54] = 16'b11111_110011_00111;
end_screen[57][55] = 16'b11111_110011_00111;
end_screen[57][56] = 16'b11111_110011_00111;
end_screen[57][57] = 16'b11111_110011_00111;
end_screen[57][58] = 16'b10001_101010_11100;
end_screen[57][59] = 16'b10001_101010_11100;
end_screen[57][60] = 16'b10001_101010_11100;
end_screen[57][61] = 16'b10001_101010_11100;
end_screen[57][62] = 16'b10001_101010_11100;
end_screen[57][63] = 16'b10001_101010_11100;
end_screen[57][64] = 16'b10001_101010_11100;
end_screen[57][65] = 16'b10001_101010_11100;
end_screen[57][66] = 16'b10001_101010_11100;
end_screen[57][67] = 16'b10001_101010_11100;
end_screen[57][68] = 16'b10001_101010_11100;
end_screen[57][69] = 16'b10001_101010_11100;
end_screen[57][70] = 16'b10001_101010_11100;
end_screen[57][71] = 16'b10001_101010_11100;
end_screen[57][72] = 16'b10001_101010_11100;
end_screen[57][73] = 16'b10001_101010_11011;
end_screen[57][74] = 16'b10110_101000_10000;
end_screen[57][75] = 16'b10111_101000_10000;
end_screen[57][76] = 16'b10111_101000_10000;
end_screen[57][77] = 16'b10111_101001_10000;
end_screen[57][78] = 16'b10111_101001_10000;
end_screen[57][79] = 16'b10111_101001_10000;
end_screen[57][80] = 16'b10111_101001_10001;
end_screen[57][81] = 16'b10111_101001_10001;
end_screen[57][82] = 16'b10111_101001_10000;
end_screen[57][83] = 16'b10111_101001_10000;
end_screen[57][84] = 16'b10001_101010_11100;
end_screen[57][85] = 16'b10001_101010_11100;
end_screen[57][86] = 16'b10001_101010_11100;
end_screen[57][87] = 16'b10001_101010_11100;
end_screen[57][88] = 16'b10001_101010_11100;
end_screen[57][89] = 16'b10001_101010_11100;
end_screen[57][90] = 16'b10001_101010_11100;
end_screen[57][91] = 16'b10001_101010_11100;
end_screen[57][92] = 16'b10001_101010_11100;
end_screen[57][93] = 16'b10001_101010_11100;
end_screen[57][94] = 16'b10001_101010_11100;
end_screen[57][95] = 16'b10001_101010_11100;
end_screen[58][0] = 16'b10001_101010_11100;
end_screen[58][1] = 16'b10001_101010_11100;
end_screen[58][2] = 16'b10001_101010_11100;
end_screen[58][3] = 16'b10001_101010_11100;
end_screen[58][4] = 16'b10001_101010_11100;
end_screen[58][5] = 16'b10001_101010_11100;
end_screen[58][6] = 16'b10001_101010_11100;
end_screen[58][7] = 16'b10001_101010_11100;
end_screen[58][8] = 16'b10001_101010_11100;
end_screen[58][9] = 16'b10001_101010_11100;
end_screen[58][10] = 16'b10010_101001_11010;
end_screen[58][11] = 16'b10100_101001_10101;
end_screen[58][12] = 16'b10101_101011_10110;
end_screen[58][13] = 16'b10101_101011_10110;
end_screen[58][14] = 16'b11010_101011_01101;
end_screen[58][15] = 16'b11010_101010_01101;
end_screen[58][16] = 16'b11010_101100_01110;
end_screen[58][17] = 16'b11011_101110_01111;
end_screen[58][18] = 16'b11011_101101_01111;
end_screen[58][19] = 16'b11011_101110_01111;
end_screen[58][20] = 16'b11100_110000_10000;
end_screen[58][21] = 16'b11011_101110_01111;
end_screen[58][22] = 16'b10110_101100_10101;
end_screen[58][23] = 16'b10101_101100_10111;
end_screen[58][24] = 16'b10110_101101_10111;
end_screen[58][25] = 16'b10101_101011_10110;
end_screen[58][26] = 16'b10011_101010_11001;
end_screen[58][27] = 16'b10001_101010_11100;
end_screen[58][28] = 16'b10001_101010_11100;
end_screen[58][29] = 16'b10001_101010_11100;
end_screen[58][30] = 16'b10001_101010_11100;
end_screen[58][31] = 16'b10001_101010_11100;
end_screen[58][32] = 16'b10001_101010_11100;
end_screen[58][33] = 16'b10001_101010_11100;
end_screen[58][34] = 16'b10001_101010_11100;
end_screen[58][35] = 16'b10001_101010_11100;
end_screen[58][36] = 16'b10001_101010_11100;
end_screen[58][37] = 16'b10001_101010_11100;
end_screen[58][38] = 16'b10001_101010_11100;
end_screen[58][39] = 16'b11111_110011_00111;
end_screen[58][40] = 16'b11111_110011_00111;
end_screen[58][41] = 16'b11111_110011_00111;
end_screen[58][42] = 16'b11111_110011_00111;
end_screen[58][43] = 16'b10001_101010_11100;
end_screen[58][44] = 16'b10001_101010_11100;
end_screen[58][45] = 16'b10001_101010_11100;
end_screen[58][46] = 16'b10001_101010_11100;
end_screen[58][47] = 16'b10001_101010_11100;
end_screen[58][48] = 16'b10001_101010_11100;
end_screen[58][49] = 16'b10001_101010_11100;
end_screen[58][50] = 16'b10001_101010_11100;
end_screen[58][51] = 16'b10001_101010_11100;
end_screen[58][52] = 16'b10001_101010_11100;
end_screen[58][53] = 16'b10001_101010_11100;
end_screen[58][54] = 16'b11111_110011_00111;
end_screen[58][55] = 16'b11111_110011_00111;
end_screen[58][56] = 16'b11111_110011_00111;
end_screen[58][57] = 16'b11111_110011_00111;
end_screen[58][58] = 16'b10001_101010_11100;
end_screen[58][59] = 16'b10001_101010_11100;
end_screen[58][60] = 16'b10001_101010_11100;
end_screen[58][61] = 16'b10001_101010_11100;
end_screen[58][62] = 16'b10001_101010_11100;
end_screen[58][63] = 16'b10001_101010_11100;
end_screen[58][64] = 16'b10001_101010_11100;
end_screen[58][65] = 16'b10001_101010_11100;
end_screen[58][66] = 16'b10001_101010_11100;
end_screen[58][67] = 16'b10001_101010_11100;
end_screen[58][68] = 16'b10001_101010_11100;
end_screen[58][69] = 16'b10001_101010_11100;
end_screen[58][70] = 16'b10001_101010_11100;
end_screen[58][71] = 16'b10001_101010_11100;
end_screen[58][72] = 16'b10001_101010_11100;
end_screen[58][73] = 16'b10001_101010_11100;
end_screen[58][74] = 16'b10001_101010_11100;
end_screen[58][75] = 16'b10001_101010_11100;
end_screen[58][76] = 16'b10001_101010_11100;
end_screen[58][77] = 16'b10001_101010_11100;
end_screen[58][78] = 16'b10001_101010_11100;
end_screen[58][79] = 16'b10001_101010_11100;
end_screen[58][80] = 16'b10001_101010_11100;
end_screen[58][81] = 16'b10001_101010_11100;
end_screen[58][82] = 16'b10001_101010_11100;
end_screen[58][83] = 16'b10001_101010_11100;
end_screen[58][84] = 16'b10001_101010_11100;
end_screen[58][85] = 16'b10001_101010_11100;
end_screen[58][86] = 16'b10001_101010_11100;
end_screen[58][87] = 16'b10001_101010_11100;
end_screen[58][88] = 16'b10001_101010_11100;
end_screen[58][89] = 16'b10001_101010_11100;
end_screen[58][90] = 16'b10001_101010_11100;
end_screen[58][91] = 16'b10001_101010_11100;
end_screen[58][92] = 16'b10001_101010_11100;
end_screen[58][93] = 16'b10001_101010_11100;
end_screen[58][94] = 16'b10001_101010_11100;
end_screen[58][95] = 16'b10001_101010_11100;
end_screen[59][0] = 16'b10001_101010_11100;
end_screen[59][1] = 16'b10001_101010_11100;
end_screen[59][2] = 16'b10001_101010_11100;
end_screen[59][3] = 16'b10001_101010_11100;
end_screen[59][4] = 16'b10001_101010_11100;
end_screen[59][5] = 16'b10001_101010_11100;
end_screen[59][6] = 16'b10001_101010_11100;
end_screen[59][7] = 16'b10001_101010_11100;
end_screen[59][8] = 16'b10001_101010_11100;
end_screen[59][9] = 16'b10001_101010_11100;
end_screen[59][10] = 16'b10001_101010_11100;
end_screen[59][11] = 16'b10001_101010_11100;
end_screen[59][12] = 16'b10001_101010_11100;
end_screen[59][13] = 16'b10001_101010_11100;
end_screen[59][14] = 16'b10100_101001_10101;
end_screen[59][15] = 16'b10101_101001_10100;
end_screen[59][16] = 16'b10101_101010_10100;
end_screen[59][17] = 16'b10110_101010_10100;
end_screen[59][18] = 16'b10110_101010_10100;
end_screen[59][19] = 16'b10110_101011_10101;
end_screen[59][20] = 16'b10111_101101_10110;
end_screen[59][21] = 16'b10110_101010_10100;
end_screen[59][22] = 16'b10001_101010_11100;
end_screen[59][23] = 16'b10001_101010_11100;
end_screen[59][24] = 16'b10001_101010_11100;
end_screen[59][25] = 16'b10001_101010_11100;
end_screen[59][26] = 16'b10001_101010_11100;
end_screen[59][27] = 16'b10001_101010_11100;
end_screen[59][28] = 16'b10001_101010_11100;
end_screen[59][29] = 16'b10001_101010_11100;
end_screen[59][30] = 16'b10001_101010_11100;
end_screen[59][31] = 16'b10001_101010_11100;
end_screen[59][32] = 16'b10001_101010_11100;
end_screen[59][33] = 16'b10001_101010_11100;
end_screen[59][34] = 16'b10001_101010_11100;
end_screen[59][35] = 16'b10001_101010_11100;
end_screen[59][36] = 16'b10001_101010_11100;
end_screen[59][37] = 16'b10001_101010_11100;
end_screen[59][38] = 16'b10001_101010_11100;
end_screen[59][39] = 16'b11111_110011_00111;
end_screen[59][40] = 16'b11111_110011_00111;
end_screen[59][41] = 16'b11111_110011_00111;
end_screen[59][42] = 16'b11111_110011_00111;
end_screen[59][43] = 16'b10001_101010_11100;
end_screen[59][44] = 16'b10001_101010_11100;
end_screen[59][45] = 16'b10001_101010_11100;
end_screen[59][46] = 16'b10001_101010_11100;
end_screen[59][47] = 16'b10001_101010_11100;
end_screen[59][48] = 16'b10001_101010_11100;
end_screen[59][49] = 16'b10001_101010_11100;
end_screen[59][50] = 16'b10001_101010_11100;
end_screen[59][51] = 16'b10001_101010_11100;
end_screen[59][52] = 16'b10001_101010_11100;
end_screen[59][53] = 16'b10001_101010_11100;
end_screen[59][54] = 16'b11111_110011_00111;
end_screen[59][55] = 16'b11111_110011_00111;
end_screen[59][56] = 16'b11111_110011_00111;
end_screen[59][57] = 16'b11111_110011_00111;
end_screen[59][58] = 16'b10001_101010_11100;
end_screen[59][59] = 16'b10001_101010_11100;
end_screen[59][60] = 16'b10001_101010_11100;
end_screen[59][61] = 16'b10001_101010_11100;
end_screen[59][62] = 16'b10001_101010_11100;
end_screen[59][63] = 16'b10001_101010_11100;
end_screen[59][64] = 16'b10001_101010_11100;
end_screen[59][65] = 16'b10001_101010_11100;
end_screen[59][66] = 16'b10001_101010_11100;
end_screen[59][67] = 16'b10001_101010_11100;
end_screen[59][68] = 16'b10001_101010_11100;
end_screen[59][69] = 16'b10001_101010_11100;
end_screen[59][70] = 16'b10001_101010_11100;
end_screen[59][71] = 16'b10001_101010_11100;
end_screen[59][72] = 16'b10001_101010_11100;
end_screen[59][73] = 16'b10001_101010_11100;
end_screen[59][74] = 16'b10001_101010_11100;
end_screen[59][75] = 16'b10001_101010_11100;
end_screen[59][76] = 16'b10001_101010_11100;
end_screen[59][77] = 16'b10001_101010_11100;
end_screen[59][78] = 16'b10001_101010_11100;
end_screen[59][79] = 16'b10001_101010_11100;
end_screen[59][80] = 16'b10001_101010_11100;
end_screen[59][81] = 16'b10001_101010_11100;
end_screen[59][82] = 16'b10001_101010_11100;
end_screen[59][83] = 16'b10001_101010_11100;
end_screen[59][84] = 16'b10001_101010_11100;
end_screen[59][85] = 16'b10001_101010_11100;
end_screen[59][86] = 16'b10001_101010_11100;
end_screen[59][87] = 16'b10001_101010_11100;
end_screen[59][88] = 16'b10001_101010_11100;
end_screen[59][89] = 16'b10001_101010_11100;
end_screen[59][90] = 16'b10001_101010_11100;
end_screen[59][91] = 16'b10001_101010_11100;
end_screen[59][92] = 16'b10001_101010_11100;
end_screen[59][93] = 16'b10001_101010_11100;
end_screen[59][94] = 16'b10001_101010_11100;
end_screen[59][95] = 16'b10001_101010_11100;
end_screen[60][0] = 16'b10001_101010_11100;
end_screen[60][1] = 16'b10001_101010_11100;
end_screen[60][2] = 16'b10001_101010_11100;
end_screen[60][3] = 16'b10001_101010_11100;
end_screen[60][4] = 16'b10001_101010_11100;
end_screen[60][5] = 16'b10001_101010_11100;
end_screen[60][6] = 16'b10001_101010_11100;
end_screen[60][7] = 16'b10001_101010_11100;
end_screen[60][8] = 16'b10001_101010_11100;
end_screen[60][9] = 16'b10001_101010_11100;
end_screen[60][10] = 16'b10001_101010_11100;
end_screen[60][11] = 16'b10001_101010_11100;
end_screen[60][12] = 16'b10001_101010_11100;
end_screen[60][13] = 16'b10001_101010_11100;
end_screen[60][14] = 16'b10001_101010_11100;
end_screen[60][15] = 16'b10001_101010_11100;
end_screen[60][16] = 16'b10001_101010_11100;
end_screen[60][17] = 16'b10001_101010_11100;
end_screen[60][18] = 16'b10001_101010_11100;
end_screen[60][19] = 16'b10001_101010_11100;
end_screen[60][20] = 16'b10001_101010_11100;
end_screen[60][21] = 16'b10001_101010_11100;
end_screen[60][22] = 16'b10001_101010_11100;
end_screen[60][23] = 16'b10001_101010_11100;
end_screen[60][24] = 16'b10001_101010_11100;
end_screen[60][25] = 16'b10001_101010_11100;
end_screen[60][26] = 16'b10001_101010_11100;
end_screen[60][27] = 16'b10001_101010_11100;
end_screen[60][28] = 16'b10001_101010_11100;
end_screen[60][29] = 16'b10001_101010_11100;
end_screen[60][30] = 16'b10001_101010_11100;
end_screen[60][31] = 16'b10001_101010_11100;
end_screen[60][32] = 16'b10001_101010_11100;
end_screen[60][33] = 16'b10001_101010_11100;
end_screen[60][34] = 16'b10001_101010_11100;
end_screen[60][35] = 16'b10001_101010_11100;
end_screen[60][36] = 16'b10001_101010_11100;
end_screen[60][37] = 16'b10001_101010_11100;
end_screen[60][38] = 16'b10001_101010_11100;
end_screen[60][39] = 16'b10001_101010_11100;
end_screen[60][40] = 16'b10001_101010_11100;
end_screen[60][41] = 16'b10001_101010_11100;
end_screen[60][42] = 16'b10001_101010_11100;
end_screen[60][43] = 16'b10001_101010_11100;
end_screen[60][44] = 16'b10001_101010_11100;
end_screen[60][45] = 16'b10001_101010_11100;
end_screen[60][46] = 16'b10001_101010_11100;
end_screen[60][47] = 16'b10001_101010_11100;
end_screen[60][48] = 16'b10001_101010_11100;
end_screen[60][49] = 16'b10001_101010_11100;
end_screen[60][50] = 16'b10001_101010_11100;
end_screen[60][51] = 16'b10001_101010_11100;
end_screen[60][52] = 16'b10001_101010_11100;
end_screen[60][53] = 16'b10001_101010_11100;
end_screen[60][54] = 16'b10001_101010_11100;
end_screen[60][55] = 16'b10001_101010_11100;
end_screen[60][56] = 16'b10001_101010_11100;
end_screen[60][57] = 16'b10001_101010_11100;
end_screen[60][58] = 16'b10001_101010_11100;
end_screen[60][59] = 16'b10001_101010_11100;
end_screen[60][60] = 16'b10001_101010_11100;
end_screen[60][61] = 16'b10001_101010_11100;
end_screen[60][62] = 16'b10001_101010_11100;
end_screen[60][63] = 16'b10001_101010_11100;
end_screen[60][64] = 16'b10001_101010_11100;
end_screen[60][65] = 16'b10001_101010_11100;
end_screen[60][66] = 16'b10001_101010_11100;
end_screen[60][67] = 16'b10001_101010_11100;
end_screen[60][68] = 16'b10001_101010_11100;
end_screen[60][69] = 16'b10001_101010_11100;
end_screen[60][70] = 16'b10001_101010_11100;
end_screen[60][71] = 16'b10001_101010_11100;
end_screen[60][72] = 16'b10001_101010_11100;
end_screen[60][73] = 16'b10001_101010_11100;
end_screen[60][74] = 16'b10001_101010_11100;
end_screen[60][75] = 16'b10001_101010_11100;
end_screen[60][76] = 16'b10001_101010_11100;
end_screen[60][77] = 16'b10001_101010_11100;
end_screen[60][78] = 16'b10001_101010_11100;
end_screen[60][79] = 16'b10001_101010_11100;
end_screen[60][80] = 16'b10001_101010_11100;
end_screen[60][81] = 16'b10001_101010_11100;
end_screen[60][82] = 16'b10001_101010_11100;
end_screen[60][83] = 16'b10001_101010_11100;
end_screen[60][84] = 16'b10001_101010_11100;
end_screen[60][85] = 16'b10001_101010_11100;
end_screen[60][86] = 16'b10001_101010_11100;
end_screen[60][87] = 16'b10001_101010_11100;
end_screen[60][88] = 16'b10001_101010_11100;
end_screen[60][89] = 16'b10001_101010_11100;
end_screen[60][90] = 16'b10001_101010_11100;
end_screen[60][91] = 16'b10001_101010_11100;
end_screen[60][92] = 16'b10001_101010_11100;
end_screen[60][93] = 16'b10001_101010_11100;
end_screen[60][94] = 16'b10001_101010_11100;
end_screen[60][95] = 16'b10001_101010_11100;
end_screen[61][0] = 16'b10001_101010_11100;
end_screen[61][1] = 16'b10001_101010_11100;
end_screen[61][2] = 16'b10001_101010_11100;
end_screen[61][3] = 16'b10001_101010_11100;
end_screen[61][4] = 16'b10001_101010_11100;
end_screen[61][5] = 16'b10001_101010_11100;
end_screen[61][6] = 16'b10001_101010_11100;
end_screen[61][7] = 16'b10001_101010_11100;
end_screen[61][8] = 16'b10001_101010_11100;
end_screen[61][9] = 16'b10001_101010_11100;
end_screen[61][10] = 16'b10001_101010_11100;
end_screen[61][11] = 16'b10001_101010_11100;
end_screen[61][12] = 16'b10001_101010_11100;
end_screen[61][13] = 16'b10001_101010_11100;
end_screen[61][14] = 16'b10001_101010_11100;
end_screen[61][15] = 16'b10001_101010_11100;
end_screen[61][16] = 16'b10001_101010_11100;
end_screen[61][17] = 16'b10001_101010_11100;
end_screen[61][18] = 16'b10001_101010_11100;
end_screen[61][19] = 16'b10001_101010_11100;
end_screen[61][20] = 16'b10001_101010_11100;
end_screen[61][21] = 16'b10001_101010_11100;
end_screen[61][22] = 16'b10001_101010_11100;
end_screen[61][23] = 16'b10001_101010_11100;
end_screen[61][24] = 16'b10001_101010_11100;
end_screen[61][25] = 16'b10001_101010_11100;
end_screen[61][26] = 16'b10001_101010_11100;
end_screen[61][27] = 16'b10001_101010_11100;
end_screen[61][28] = 16'b10001_101010_11100;
end_screen[61][29] = 16'b10001_101010_11100;
end_screen[61][30] = 16'b10001_101010_11100;
end_screen[61][31] = 16'b10001_101010_11100;
end_screen[61][32] = 16'b10001_101010_11100;
end_screen[61][33] = 16'b10001_101010_11100;
end_screen[61][34] = 16'b10001_101010_11100;
end_screen[61][35] = 16'b10001_101010_11100;
end_screen[61][36] = 16'b10001_101010_11100;
end_screen[61][37] = 16'b10001_101010_11100;
end_screen[61][38] = 16'b10001_101010_11100;
end_screen[61][39] = 16'b10001_101010_11100;
end_screen[61][40] = 16'b10001_101010_11100;
end_screen[61][41] = 16'b10001_101010_11100;
end_screen[61][42] = 16'b10001_101010_11100;
end_screen[61][43] = 16'b10001_101010_11100;
end_screen[61][44] = 16'b10001_101010_11100;
end_screen[61][45] = 16'b10001_101010_11100;
end_screen[61][46] = 16'b10001_101010_11100;
end_screen[61][47] = 16'b10001_101010_11100;
end_screen[61][48] = 16'b10001_101010_11100;
end_screen[61][49] = 16'b10001_101010_11100;
end_screen[61][50] = 16'b10001_101010_11100;
end_screen[61][51] = 16'b10001_101010_11100;
end_screen[61][52] = 16'b10001_101010_11100;
end_screen[61][53] = 16'b10001_101010_11100;
end_screen[61][54] = 16'b10001_101010_11100;
end_screen[61][55] = 16'b10001_101010_11100;
end_screen[61][56] = 16'b10001_101010_11100;
end_screen[61][57] = 16'b10001_101010_11100;
end_screen[61][58] = 16'b10001_101010_11100;
end_screen[61][59] = 16'b10001_101010_11100;
end_screen[61][60] = 16'b10001_101010_11100;
end_screen[61][61] = 16'b10001_101010_11100;
end_screen[61][62] = 16'b10001_101010_11100;
end_screen[61][63] = 16'b10001_101010_11100;
end_screen[61][64] = 16'b10001_101010_11100;
end_screen[61][65] = 16'b10001_101010_11100;
end_screen[61][66] = 16'b10001_101010_11100;
end_screen[61][67] = 16'b10001_101010_11100;
end_screen[61][68] = 16'b10001_101010_11100;
end_screen[61][69] = 16'b10001_101010_11100;
end_screen[61][70] = 16'b10001_101010_11100;
end_screen[61][71] = 16'b10001_101010_11100;
end_screen[61][72] = 16'b10001_101010_11100;
end_screen[61][73] = 16'b10001_101010_11100;
end_screen[61][74] = 16'b10001_101010_11100;
end_screen[61][75] = 16'b10001_101010_11100;
end_screen[61][76] = 16'b10001_101010_11100;
end_screen[61][77] = 16'b10001_101010_11100;
end_screen[61][78] = 16'b10001_101010_11100;
end_screen[61][79] = 16'b10001_101010_11100;
end_screen[61][80] = 16'b10001_101010_11100;
end_screen[61][81] = 16'b10001_101010_11100;
end_screen[61][82] = 16'b10001_101010_11100;
end_screen[61][83] = 16'b10001_101010_11100;
end_screen[61][84] = 16'b10001_101010_11100;
end_screen[61][85] = 16'b10001_101010_11100;
end_screen[61][86] = 16'b10001_101010_11100;
end_screen[61][87] = 16'b10001_101010_11100;
end_screen[61][88] = 16'b10001_101010_11100;
end_screen[61][89] = 16'b10001_101010_11100;
end_screen[61][90] = 16'b10001_101010_11100;
end_screen[61][91] = 16'b10001_101010_11100;
end_screen[61][92] = 16'b10001_101010_11100;
end_screen[61][93] = 16'b10001_101010_11100;
end_screen[61][94] = 16'b10001_101010_11100;
end_screen[61][95] = 16'b10001_101010_11100;
end_screen[62][0] = 16'b10001_101010_11100;
end_screen[62][1] = 16'b10001_101010_11100;
end_screen[62][2] = 16'b10001_101010_11100;
end_screen[62][3] = 16'b10001_101010_11100;
end_screen[62][4] = 16'b10001_101010_11100;
end_screen[62][5] = 16'b10001_101010_11100;
end_screen[62][6] = 16'b10001_101010_11100;
end_screen[62][7] = 16'b10001_101010_11100;
end_screen[62][8] = 16'b10001_101010_11100;
end_screen[62][9] = 16'b10001_101010_11100;
end_screen[62][10] = 16'b10001_101010_11100;
end_screen[62][11] = 16'b10001_101010_11100;
end_screen[62][12] = 16'b10001_101010_11100;
end_screen[62][13] = 16'b10001_101010_11100;
end_screen[62][14] = 16'b10001_101010_11100;
end_screen[62][15] = 16'b10001_101010_11100;
end_screen[62][16] = 16'b10001_101010_11100;
end_screen[62][17] = 16'b10001_101010_11100;
end_screen[62][18] = 16'b10001_101010_11100;
end_screen[62][19] = 16'b10001_101010_11100;
end_screen[62][20] = 16'b10001_101010_11100;
end_screen[62][21] = 16'b10001_101010_11100;
end_screen[62][22] = 16'b10001_101010_11100;
end_screen[62][23] = 16'b10001_101010_11100;
end_screen[62][24] = 16'b10001_101010_11100;
end_screen[62][25] = 16'b10001_101010_11100;
end_screen[62][26] = 16'b10001_101010_11100;
end_screen[62][27] = 16'b10001_101010_11100;
end_screen[62][28] = 16'b10001_101010_11100;
end_screen[62][29] = 16'b10001_101010_11100;
end_screen[62][30] = 16'b10001_101010_11100;
end_screen[62][31] = 16'b10001_101010_11100;
end_screen[62][32] = 16'b10001_101010_11100;
end_screen[62][33] = 16'b10001_101010_11100;
end_screen[62][34] = 16'b10001_101010_11100;
end_screen[62][35] = 16'b10001_101010_11100;
end_screen[62][36] = 16'b10001_101010_11100;
end_screen[62][37] = 16'b10001_101010_11100;
end_screen[62][38] = 16'b10001_101010_11100;
end_screen[62][39] = 16'b10001_101010_11100;
end_screen[62][40] = 16'b10001_101010_11100;
end_screen[62][41] = 16'b10001_101010_11100;
end_screen[62][42] = 16'b10001_101010_11100;
end_screen[62][43] = 16'b10001_101010_11100;
end_screen[62][44] = 16'b10001_101010_11100;
end_screen[62][45] = 16'b10001_101010_11100;
end_screen[62][46] = 16'b10001_101010_11100;
end_screen[62][47] = 16'b10001_101010_11100;
end_screen[62][48] = 16'b10001_101010_11100;
end_screen[62][49] = 16'b10001_101010_11100;
end_screen[62][50] = 16'b10001_101010_11100;
end_screen[62][51] = 16'b10001_101010_11100;
end_screen[62][52] = 16'b10001_101010_11100;
end_screen[62][53] = 16'b10001_101010_11100;
end_screen[62][54] = 16'b10001_101010_11100;
end_screen[62][55] = 16'b10001_101010_11100;
end_screen[62][56] = 16'b10001_101010_11100;
end_screen[62][57] = 16'b10001_101010_11100;
end_screen[62][58] = 16'b10001_101010_11100;
end_screen[62][59] = 16'b10001_101010_11100;
end_screen[62][60] = 16'b10001_101010_11100;
end_screen[62][61] = 16'b10001_101010_11100;
end_screen[62][62] = 16'b10001_101010_11100;
end_screen[62][63] = 16'b10001_101010_11100;
end_screen[62][64] = 16'b10001_101010_11100;
end_screen[62][65] = 16'b10001_101010_11100;
end_screen[62][66] = 16'b10001_101010_11100;
end_screen[62][67] = 16'b10001_101010_11100;
end_screen[62][68] = 16'b10001_101010_11100;
end_screen[62][69] = 16'b10001_101010_11100;
end_screen[62][70] = 16'b10001_101010_11100;
end_screen[62][71] = 16'b10001_101010_11100;
end_screen[62][72] = 16'b10001_101010_11100;
end_screen[62][73] = 16'b10001_101010_11100;
end_screen[62][74] = 16'b10001_101010_11100;
end_screen[62][75] = 16'b10001_101010_11100;
end_screen[62][76] = 16'b10001_101010_11100;
end_screen[62][77] = 16'b10001_101010_11100;
end_screen[62][78] = 16'b10001_101010_11100;
end_screen[62][79] = 16'b10001_101010_11100;
end_screen[62][80] = 16'b10001_101010_11100;
end_screen[62][81] = 16'b10001_101010_11100;
end_screen[62][82] = 16'b10001_101010_11100;
end_screen[62][83] = 16'b10001_101010_11100;
end_screen[62][84] = 16'b10001_101010_11100;
end_screen[62][85] = 16'b10001_101010_11100;
end_screen[62][86] = 16'b10001_101010_11100;
end_screen[62][87] = 16'b10001_101010_11100;
end_screen[62][88] = 16'b10001_101010_11100;
end_screen[62][89] = 16'b10001_101010_11100;
end_screen[62][90] = 16'b10001_101010_11100;
end_screen[62][91] = 16'b10001_101010_11100;
end_screen[62][92] = 16'b10001_101010_11100;
end_screen[62][93] = 16'b10001_101010_11100;
end_screen[62][94] = 16'b10001_101010_11100;
end_screen[62][95] = 16'b10001_101010_11100;
end_screen[63][0] = 16'b10001_101010_11100;
end_screen[63][1] = 16'b10001_101010_11100;
end_screen[63][2] = 16'b10001_101010_11100;
end_screen[63][3] = 16'b10001_101010_11100;
end_screen[63][4] = 16'b10001_101010_11100;
end_screen[63][5] = 16'b10001_101010_11100;
end_screen[63][6] = 16'b10001_101010_11100;
end_screen[63][7] = 16'b10001_101010_11100;
end_screen[63][8] = 16'b10001_101010_11100;
end_screen[63][9] = 16'b10001_101010_11100;
end_screen[63][10] = 16'b10001_101010_11100;
end_screen[63][11] = 16'b10001_101010_11100;
end_screen[63][12] = 16'b10001_101010_11100;
end_screen[63][13] = 16'b10001_101010_11100;
end_screen[63][14] = 16'b10001_101010_11100;
end_screen[63][15] = 16'b10001_101010_11100;
end_screen[63][16] = 16'b10001_101010_11100;
end_screen[63][17] = 16'b10001_101010_11100;
end_screen[63][18] = 16'b10001_101010_11100;
end_screen[63][19] = 16'b10001_101010_11100;
end_screen[63][20] = 16'b10001_101010_11100;
end_screen[63][21] = 16'b10001_101010_11100;
end_screen[63][22] = 16'b10001_101010_11100;
end_screen[63][23] = 16'b10001_101010_11100;
end_screen[63][24] = 16'b10001_101010_11100;
end_screen[63][25] = 16'b10001_101010_11100;
end_screen[63][26] = 16'b10001_101010_11100;
end_screen[63][27] = 16'b10001_101010_11100;
end_screen[63][28] = 16'b10001_101010_11100;
end_screen[63][29] = 16'b10001_101010_11100;
end_screen[63][30] = 16'b10001_101010_11100;
end_screen[63][31] = 16'b10001_101010_11100;
end_screen[63][32] = 16'b10001_101010_11100;
end_screen[63][33] = 16'b10001_101010_11100;
end_screen[63][34] = 16'b10001_101010_11100;
end_screen[63][35] = 16'b10001_101010_11100;
end_screen[63][36] = 16'b10001_101010_11100;
end_screen[63][37] = 16'b10001_101010_11100;
end_screen[63][38] = 16'b10001_101010_11100;
end_screen[63][39] = 16'b10001_101010_11100;
end_screen[63][40] = 16'b10001_101010_11100;
end_screen[63][41] = 16'b10001_101010_11100;
end_screen[63][42] = 16'b10001_101010_11100;
end_screen[63][43] = 16'b10001_101010_11100;
end_screen[63][44] = 16'b10001_101010_11100;
end_screen[63][45] = 16'b10001_101010_11100;
end_screen[63][46] = 16'b10001_101010_11100;
end_screen[63][47] = 16'b10001_101010_11100;
end_screen[63][48] = 16'b10001_101010_11100;
end_screen[63][49] = 16'b10001_101010_11100;
end_screen[63][50] = 16'b10001_101010_11100;
end_screen[63][51] = 16'b10001_101010_11100;
end_screen[63][52] = 16'b10001_101010_11100;
end_screen[63][53] = 16'b10001_101010_11100;
end_screen[63][54] = 16'b10001_101010_11100;
end_screen[63][55] = 16'b10001_101010_11100;
end_screen[63][56] = 16'b10001_101010_11100;
end_screen[63][57] = 16'b10001_101010_11100;
end_screen[63][58] = 16'b10001_101010_11100;
end_screen[63][59] = 16'b10001_101010_11100;
end_screen[63][60] = 16'b10001_101010_11100;
end_screen[63][61] = 16'b10001_101010_11100;
end_screen[63][62] = 16'b10001_101010_11100;
end_screen[63][63] = 16'b10001_101010_11100;
end_screen[63][64] = 16'b10001_101010_11100;
end_screen[63][65] = 16'b10001_101010_11100;
end_screen[63][66] = 16'b10001_101010_11100;
end_screen[63][67] = 16'b10001_101010_11100;
end_screen[63][68] = 16'b10001_101010_11100;
end_screen[63][69] = 16'b10001_101010_11100;
end_screen[63][70] = 16'b10001_101010_11100;
end_screen[63][71] = 16'b10001_101010_11100;
end_screen[63][72] = 16'b10001_101010_11100;
end_screen[63][73] = 16'b10001_101010_11100;
end_screen[63][74] = 16'b10001_101010_11100;
end_screen[63][75] = 16'b10001_101010_11100;
end_screen[63][76] = 16'b10001_101010_11100;
end_screen[63][77] = 16'b10001_101010_11100;
end_screen[63][78] = 16'b10001_101010_11100;
end_screen[63][79] = 16'b10001_101010_11100;
end_screen[63][80] = 16'b10001_101010_11100;
end_screen[63][81] = 16'b10001_101010_11100;
end_screen[63][82] = 16'b10001_101010_11100;
end_screen[63][83] = 16'b10001_101010_11100;
end_screen[63][84] = 16'b10001_101010_11100;
end_screen[63][85] = 16'b10001_101010_11100;
end_screen[63][86] = 16'b10001_101010_11100;
end_screen[63][87] = 16'b10001_101010_11100;
end_screen[63][88] = 16'b10001_101010_11100;
end_screen[63][89] = 16'b10001_101010_11100;
end_screen[63][90] = 16'b10001_101010_11100;
end_screen[63][91] = 16'b10001_101010_11100;
end_screen[63][92] = 16'b10001_101010_11100;
end_screen[63][93] = 16'b10001_101010_11100;
end_screen[63][94] = 16'b10001_101010_11100;
end_screen[63][95] = 16'b10001_101010_11100;

end

always @ (posedge basys_clk) begin
    oled_data <= end_screen[y][x];
end

endmodule
