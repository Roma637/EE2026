`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09.04.2025 11:10:35
// Design Name: 
// Module Name: draw_ingredients
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module draw_ingredients#(
    parameter ONION_TOP_LEFT_X = 2,
    parameter ONION_TOP_LEFT_Y = 2,
    parameter TOMATO_TOP_LEFT_X = 2,
    parameter TOMATO_TOP_LEFT_Y = 47,
    parameter CHICKEN_TOP_LEFT_X = 30,
    parameter CHICKEN_TOP_LEFT_Y = 47,
    parameter RICE_TOP_LEFT_X = 51,
    parameter RICE_TOP_LEFT_Y = 2
)(
    input clk_25MHz,
    input [7:0] x,
    input [6:0] y,
    output reg [15:0] oled_data 
    );
    
    reg [15:0] onion [0:14] [0:14];
    reg [15:0] rice [0:14] [0:14];
    reg [15:0] tomato [0:14] [0:14];
    reg [15:0] chicken [0:14] [0:14];
    
    // set x,y of top left hand corner of zones here!!
    
    reg [7:0] onion_x_offset = 0 ;
    reg [6:0] onion_y_offset = 0 ;
    
    reg [7:0] rice_x_offset = 20 ;
    reg [6:0] rice_y_offset = 0 ;
    
    reg [7:0] chicken_x_offset = 0 ;
    reg [6:0] chicken_y_offset = 20 ;
    
    reg [7:0] tomato_x_offset = 20 ;
    reg [6:0] tomato_y_offset = 20 ;
    
    initial begin
        onion[0][0] = 16'b11001_100101_11111;
        onion[0][1] = 16'b11001_100101_11111;
        onion[0][2] = 16'b11001_100101_11111;
        onion[0][3] = 16'b11001_100101_11111;
        onion[0][4] = 16'b11001_100101_11111;
        onion[0][5] = 16'b11001_100101_11111;
        onion[0][6] = 16'b11001_100101_11111;
        onion[0][7] = 16'b11001_100101_11111;
        onion[0][8] = 16'b11001_100101_11111;
        onion[0][9] = 16'b11001_100101_11111;
        onion[0][10] = 16'b11001_100101_11111;
        onion[0][11] = 16'b11001_100101_11111;
        onion[0][12] = 16'b11001_100101_11111;
        onion[0][13] = 16'b11001_100101_11111;
        onion[0][14] = 16'b11001_100101_11111;
        onion[1][0] = 16'b11001_100101_11111;
        onion[1][1] = 16'b00000_000000_00000;
        onion[1][2] = 16'b00000_000000_00000;
        onion[1][3] = 16'b00000_000000_00000;
        onion[1][4] = 16'b00000_000000_00000;
        onion[1][5] = 16'b00000_000000_00000;
        onion[1][6] = 16'b00000_000000_00000;
        onion[1][7] = 16'b10100_000000_11111;
        onion[1][8] = 16'b00000_000000_00000;
        onion[1][9] = 16'b00000_000000_00000;
        onion[1][10] = 16'b00000_000000_00000;
        onion[1][11] = 16'b00000_000000_00000;
        onion[1][12] = 16'b00000_000000_00000;
        onion[1][13] = 16'b00000_000000_00000;
        onion[1][14] = 16'b11001_100101_11111;
        onion[2][0] = 16'b11001_100101_11111;
        onion[2][1] = 16'b00000_000000_00000;
        onion[2][2] = 16'b00000_000000_00000;
        onion[2][3] = 16'b00000_000000_00000;
        onion[2][4] = 16'b00000_000000_00000;
        onion[2][5] = 16'b00000_000000_00000;
        onion[2][6] = 16'b10100_000000_11111;
        onion[2][7] = 16'b11001_100101_11111;
        onion[2][8] = 16'b11001_100101_11111;
        onion[2][9] = 16'b10100_000000_11111;
        onion[2][10] = 16'b00000_000000_00000;
        onion[2][11] = 16'b00000_000000_00000;
        onion[2][12] = 16'b00000_000000_00000;
        onion[2][13] = 16'b00000_000000_00000;
        onion[2][14] = 16'b11001_100101_11111;
        onion[3][0] = 16'b11001_100101_11111;
        onion[3][1] = 16'b00000_000000_00000;
        onion[3][2] = 16'b00000_000000_00000;
        onion[3][3] = 16'b00000_000000_00000;
        onion[3][4] = 16'b00000_000000_00000;
        onion[3][5] = 16'b10100_000000_11111;
        onion[3][6] = 16'b11001_100101_11111;
        onion[3][7] = 16'b10100_000000_11111;
        onion[3][8] = 16'b10100_000000_11111;
        onion[3][9] = 16'b11001_100101_11111;
        onion[3][10] = 16'b10100_000000_11111;
        onion[3][11] = 16'b00000_000000_00000;
        onion[3][12] = 16'b00000_000000_00000;
        onion[3][13] = 16'b00000_000000_00000;
        onion[3][14] = 16'b11001_100101_11111;
        onion[4][0] = 16'b11001_100101_11111;
        onion[4][1] = 16'b00000_000000_00000;
        onion[4][2] = 16'b00000_000000_00000;
        onion[4][3] = 16'b00000_000000_00000;
        onion[4][4] = 16'b10100_000000_11111;
        onion[4][5] = 16'b11001_100101_11111;
        onion[4][6] = 16'b10100_000000_11111;
        onion[4][7] = 16'b10100_000000_11111;
        onion[4][8] = 16'b10100_000000_11111;
        onion[4][9] = 16'b10100_000000_11111;
        onion[4][10] = 16'b11001_100101_11111;
        onion[4][11] = 16'b10100_000000_11111;
        onion[4][12] = 16'b00000_000000_00000;
        onion[4][13] = 16'b00000_000000_00000;
        onion[4][14] = 16'b11001_100101_11111;
        onion[5][0] = 16'b11001_100101_11111;
        onion[5][1] = 16'b00000_000000_00000;
        onion[5][2] = 16'b00000_000000_00000;
        onion[5][3] = 16'b10100_000000_11111;
        onion[5][4] = 16'b11001_100101_11111;
        onion[5][5] = 16'b10100_000000_11111;
        onion[5][6] = 16'b10100_000000_11111;
        onion[5][7] = 16'b11001_100101_11111;
        onion[5][8] = 16'b11001_100101_11111;
        onion[5][9] = 16'b10100_000000_11111;
        onion[5][10] = 16'b10100_000000_11111;
        onion[5][11] = 16'b11001_100101_11111;
        onion[5][12] = 16'b10100_000000_11111;
        onion[5][13] = 16'b00000_000000_00000;
        onion[5][14] = 16'b11001_100101_11111;
        onion[6][0] = 16'b11001_100101_11111;
        onion[6][1] = 16'b00000_000000_00000;
        onion[6][2] = 16'b10100_000000_11111;
        onion[6][3] = 16'b11001_100101_11111;
        onion[6][4] = 16'b10100_000000_11111;
        onion[6][5] = 16'b10100_000000_11111;
        onion[6][6] = 16'b11001_100101_11111;
        onion[6][7] = 16'b10100_000000_11111;
        onion[6][8] = 16'b10100_000000_11111;
        onion[6][9] = 16'b11001_100101_11111;
        onion[6][10] = 16'b10100_000000_11111;
        onion[6][11] = 16'b10100_000000_11111;
        onion[6][12] = 16'b11001_100101_11111;
        onion[6][13] = 16'b10100_000000_11111;
        onion[6][14] = 16'b11001_100101_11111;
        onion[7][0] = 16'b11001_100101_11111;
        onion[7][1] = 16'b00000_000000_00000;
        onion[7][2] = 16'b11001_100101_11111;
        onion[7][3] = 16'b10100_000000_11111;
        onion[7][4] = 16'b10100_000000_11111;
        onion[7][5] = 16'b11001_100101_11111;
        onion[7][6] = 16'b10100_000000_11111;
        onion[7][7] = 16'b10100_000000_11111;
        onion[7][8] = 16'b11001_100101_11111;
        onion[7][9] = 16'b10100_000000_11111;
        onion[7][10] = 16'b11001_100101_11111;
        onion[7][11] = 16'b10100_000000_11111;
        onion[7][12] = 16'b11001_100101_11111;
        onion[7][13] = 16'b10100_000000_11111;
        onion[7][14] = 16'b11001_100101_11111;
        onion[8][0] = 16'b11001_100101_11111;
        onion[8][1] = 16'b10100_000000_11111;
        onion[8][2] = 16'b11001_100101_11111;
        onion[8][3] = 16'b10100_000000_11111;
        onion[8][4] = 16'b11001_100101_11111;
        onion[8][5] = 16'b10100_000000_11111;
        onion[8][6] = 16'b10100_000000_11111;
        onion[8][7] = 16'b11001_100101_11111;
        onion[8][8] = 16'b10100_000000_11111;
        onion[8][9] = 16'b10100_000000_11111;
        onion[8][10] = 16'b11001_100101_11111;
        onion[8][11] = 16'b10100_000000_11111;
        onion[8][12] = 16'b11001_100101_11111;
        onion[8][13] = 16'b10100_000000_11111;
        onion[8][14] = 16'b11001_100101_11111;
        onion[9][0] = 16'b11001_100101_11111;
        onion[9][1] = 16'b10100_000000_11111;
        onion[9][2] = 16'b11001_100101_11111;
        onion[9][3] = 16'b10100_000000_11111;
        onion[9][4] = 16'b11001_100101_11111;
        onion[9][5] = 16'b10100_000000_11111;
        onion[9][6] = 16'b10100_000000_11111;
        onion[9][7] = 16'b10100_000000_11111;
        onion[9][8] = 16'b10100_000000_11111;
        onion[9][9] = 16'b10100_000000_11111;
        onion[9][10] = 16'b11001_100101_11111;
        onion[9][11] = 16'b10100_000000_11111;
        onion[9][12] = 16'b11001_100101_11111;
        onion[9][13] = 16'b10100_000000_11111;
        onion[9][14] = 16'b11001_100101_11111;
        onion[10][0] = 16'b11001_100101_11111;
        onion[10][1] = 16'b10100_000000_11111;
        onion[10][2] = 16'b11001_100101_11111;
        onion[10][3] = 16'b10100_000000_11111;
        onion[10][4] = 16'b10100_000000_11111;
        onion[10][5] = 16'b11001_100101_11111;
        onion[10][6] = 16'b11001_100101_11111;
        onion[10][7] = 16'b11001_100101_11111;
        onion[10][8] = 16'b11001_100101_11111;
        onion[10][9] = 16'b11001_100101_11111;
        onion[10][10] = 16'b10100_000000_11111;
        onion[10][11] = 16'b10100_000000_11111;
        onion[10][12] = 16'b11001_100101_11111;
        onion[10][13] = 16'b10100_000000_11111;
        onion[10][14] = 16'b11001_100101_11111;
        onion[11][0] = 16'b11001_100101_11111;
        onion[11][1] = 16'b10100_000000_11111;
        onion[11][2] = 16'b10100_000000_11111;
        onion[11][3] = 16'b11001_100101_11111;
        onion[11][4] = 16'b10100_000000_11111;
        onion[11][5] = 16'b10100_000000_11111;
        onion[11][6] = 16'b10100_000000_11111;
        onion[11][7] = 16'b10100_000000_11111;
        onion[11][8] = 16'b10100_000000_11111;
        onion[11][9] = 16'b10100_000000_11111;
        onion[11][10] = 16'b10100_000000_11111;
        onion[11][11] = 16'b11001_100101_11111;
        onion[11][12] = 16'b10100_000000_11111;
        onion[11][13] = 16'b00000_000000_00000;
        onion[11][14] = 16'b11001_100101_11111;
        onion[12][0] = 16'b11001_100101_11111;
        onion[12][1] = 16'b00000_000000_00000;
        onion[12][2] = 16'b10100_000000_11111;
        onion[12][3] = 16'b10100_000000_11111;
        onion[12][4] = 16'b11001_100101_11111;
        onion[12][5] = 16'b11001_100101_11111;
        onion[12][6] = 16'b11001_100101_11111;
        onion[12][7] = 16'b11001_100101_11111;
        onion[12][8] = 16'b11001_100101_11111;
        onion[12][9] = 16'b11001_100101_11111;
        onion[12][10] = 16'b11001_100101_11111;
        onion[12][11] = 16'b11001_100101_11111;
        onion[12][12] = 16'b10100_000000_11111;
        onion[12][13] = 16'b00000_000000_00000;
        onion[12][14] = 16'b11001_100101_11111;
        onion[13][0] = 16'b11001_100101_11111;
        onion[13][1] = 16'b00000_000000_00000;
        onion[13][2] = 16'b00000_000000_00000;
        onion[13][3] = 16'b10100_000000_11111;
        onion[13][4] = 16'b10100_000000_11111;
        onion[13][5] = 16'b10100_000000_11111;
        onion[13][6] = 16'b10100_000000_11111;
        onion[13][7] = 16'b10100_000000_11111;
        onion[13][8] = 16'b10100_000000_11111;
        onion[13][9] = 16'b10100_000000_11111;
        onion[13][10] = 16'b10100_000000_11111;
        onion[13][11] = 16'b00000_000000_00000;
        onion[13][12] = 16'b00000_000000_00000;
        onion[13][13] = 16'b00000_000000_00000;
        onion[13][14] = 16'b11001_100101_11111;
        onion[14][0] = 16'b11001_100101_11111;
        onion[14][1] = 16'b11001_100101_11111;
        onion[14][2] = 16'b11001_100101_11111;
        onion[14][3] = 16'b11001_100101_11111;
        onion[14][4] = 16'b11001_100101_11111;
        onion[14][5] = 16'b11001_100101_11111;
        onion[14][6] = 16'b11001_100101_11111;
        onion[14][7] = 16'b11001_100101_11111;
        onion[14][8] = 16'b11001_100101_11111;
        onion[14][9] = 16'b11001_100101_11111;
        onion[14][10] = 16'b11001_100101_11111;
        onion[14][11] = 16'b11001_100101_11111;
        onion[14][12] = 16'b11001_100101_11111;
        onion[14][13] = 16'b11001_100101_11111;
        onion[14][14] = 16'b11001_100101_11111;

    
        rice[0][0] = 16'b00000_110000_11111;
        rice[0][1] = 16'b00000_110000_11111;
        rice[0][2] = 16'b00000_110000_11111;
        rice[0][3] = 16'b00000_110000_11111;
        rice[0][4] = 16'b00000_110000_11111;
        rice[0][5] = 16'b00000_110000_11111;
        rice[0][6] = 16'b00000_110000_11111;
        rice[0][7] = 16'b00000_110000_11111;
        rice[0][8] = 16'b00000_110000_11111;
        rice[0][9] = 16'b00000_110000_11111;
        rice[0][10] = 16'b00000_110000_11111;
        rice[0][11] = 16'b00000_110000_11111;
        rice[0][12] = 16'b00000_110000_11111;
        rice[0][13] = 16'b00000_110000_11111;
        rice[0][14] = 16'b00000_110000_11111;
        rice[1][0] = 16'b00000_110000_11111;
        rice[1][1] = 16'b00000_000000_00000;
        rice[1][2] = 16'b00000_000000_00000;
        rice[1][3] = 16'b00000_000000_00000;
        rice[1][4] = 16'b00000_000000_00000;
        rice[1][5] = 16'b00000_000000_00000;
        rice[1][6] = 16'b00000_000000_00000;
        rice[1][7] = 16'b00000_000000_00000;
        rice[1][8] = 16'b00000_000000_00000;
        rice[1][9] = 16'b00000_000000_00000;
        rice[1][10] = 16'b00000_000000_00000;
        rice[1][11] = 16'b00000_000000_00000;
        rice[1][12] = 16'b00000_000000_00000;
        rice[1][13] = 16'b00000_000000_00000;
        rice[1][14] = 16'b00000_110000_11111;
        rice[2][0] = 16'b00000_110000_11111;
        rice[2][1] = 16'b00000_000000_00000;
        rice[2][2] = 16'b00000_000000_00000;
        rice[2][3] = 16'b00000_000000_00000;
        rice[2][4] = 16'b00000_000000_00000;
        rice[2][5] = 16'b00000_000000_00000;
        rice[2][6] = 16'b11111_111110_11111;
        rice[2][7] = 16'b11111_111110_11111;
        rice[2][8] = 16'b11111_111110_11111;
        rice[2][9] = 16'b00000_000000_00000;
        rice[2][10] = 16'b00000_000000_00000;
        rice[2][11] = 16'b00000_000000_00000;
        rice[2][12] = 16'b00000_000000_00000;
        rice[2][13] = 16'b00000_000000_00000;
        rice[2][14] = 16'b00000_110000_11111;
        rice[3][0] = 16'b00000_110000_11111;
        rice[3][1] = 16'b00000_000000_00000;
        rice[3][2] = 16'b00000_000000_00000;
        rice[3][3] = 16'b00000_000000_00000;
        rice[3][4] = 16'b00000_000000_00000;
        rice[3][5] = 16'b11111_111111_11111;
        rice[3][6] = 16'b11111_111111_11111;
        rice[3][7] = 16'b11111_111111_11111;
        rice[3][8] = 16'b10001_100011_10001;
        rice[3][9] = 16'b11111_111111_11111;
        rice[3][10] = 16'b00000_000000_00000;
        rice[3][11] = 16'b00000_000000_00000;
        rice[3][12] = 16'b00000_000000_00000;
        rice[3][13] = 16'b00000_000000_00000;
        rice[3][14] = 16'b00000_110000_11111;
        rice[4][0] = 16'b00000_110000_11111;
        rice[4][1] = 16'b00000_000000_00000;
        rice[4][2] = 16'b00000_000000_00000;
        rice[4][3] = 16'b00000_000000_00000;
        rice[4][4] = 16'b11111_111111_11111;
        rice[4][5] = 16'b11111_111111_11111;
        rice[4][6] = 16'b10001_100011_10001;
        rice[4][7] = 16'b11111_111111_11111;
        rice[4][8] = 16'b11111_111111_11111;
        rice[4][9] = 16'b11111_111111_11111;
        rice[4][10] = 16'b11111_111111_11111;
        rice[4][11] = 16'b00000_000000_00000;
        rice[4][12] = 16'b00000_000000_00000;
        rice[4][13] = 16'b00000_000000_00000;
        rice[4][14] = 16'b00000_110000_11111;
        rice[5][0] = 16'b00000_110000_11111;
        rice[5][1] = 16'b00000_000000_00000;
        rice[5][2] = 16'b00000_000000_00000;
        rice[5][3] = 16'b11111_111111_11111;
        rice[5][4] = 16'b11111_111111_11111;
        rice[5][5] = 16'b11111_111111_11111;
        rice[5][6] = 16'b11111_111111_11111;
        rice[5][7] = 16'b11111_111111_11111;
        rice[5][8] = 16'b11111_111111_11111;
        rice[5][9] = 16'b10001_100011_10001;
        rice[5][10] = 16'b11111_111111_11111;
        rice[5][11] = 16'b11111_111111_11111;
        rice[5][12] = 16'b00000_000000_00000;
        rice[5][13] = 16'b00000_000000_00000;
        rice[5][14] = 16'b00000_110000_11111;
        rice[6][0] = 16'b00000_110000_11111;
        rice[6][1] = 16'b00000_000000_00000;
        rice[6][2] = 16'b00000_000000_00000;
        rice[6][3] = 16'b10001_100011_10001;
        rice[6][4] = 16'b11111_111111_11111;
        rice[6][5] = 16'b10001_100011_10001;
        rice[6][6] = 16'b11111_111111_11111;
        rice[6][7] = 16'b10001_100011_10001;
        rice[6][8] = 16'b11111_111111_11111;
        rice[6][9] = 16'b11111_111111_11111;
        rice[6][10] = 16'b11111_111111_11111;
        rice[6][11] = 16'b10001_100011_10001;
        rice[6][12] = 16'b00000_000000_00000;
        rice[6][13] = 16'b00000_000000_00000;
        rice[6][14] = 16'b00000_110000_11111;
        rice[7][0] = 16'b00000_110000_11111;
        rice[7][1] = 16'b00000_000000_00000;
        rice[7][2] = 16'b00000_110000_11111;
        rice[7][3] = 16'b11111_111110_11111;
        rice[7][4] = 16'b11111_111110_11111;
        rice[7][5] = 16'b11111_111110_11111;
        rice[7][6] = 16'b11111_111110_11111;
        rice[7][7] = 16'b11111_111110_11111;
        rice[7][8] = 16'b11111_111110_11111;
        rice[7][9] = 16'b10001_100011_10001;
        rice[7][10] = 16'b11111_111110_11111;
        rice[7][11] = 16'b11111_111110_11111;
        rice[7][12] = 16'b00000_110000_11111;
        rice[7][13] = 16'b00000_000000_00000;
        rice[7][14] = 16'b00000_110000_11111;
        rice[8][0] = 16'b00000_110000_11111;
        rice[8][1] = 16'b00000_000000_00000;
        rice[8][2] = 16'b00000_110000_11111;
        rice[8][3] = 16'b00000_110000_11111;
        rice[8][4] = 16'b11111_111110_11111;
        rice[8][5] = 16'b11111_111110_11111;
        rice[8][6] = 16'b10001_100011_10001;
        rice[8][7] = 16'b11111_111110_11111;
        rice[8][8] = 16'b11111_111110_11111;
        rice[8][9] = 16'b11111_111110_11111;
        rice[8][10] = 16'b11111_111110_11111;
        rice[8][11] = 16'b00000_110000_11111;
        rice[8][12] = 16'b00000_110000_11111;
        rice[8][13] = 16'b00000_000000_00000;
        rice[8][14] = 16'b00000_110000_11111;
        rice[9][0] = 16'b00000_110000_11111;
        rice[9][1] = 16'b00000_000000_00000;
        rice[9][2] = 16'b00000_110000_11111;
        rice[9][3] = 16'b00000_110000_11111;
        rice[9][4] = 16'b00000_110000_11111;
        rice[9][5] = 16'b00000_110000_11111;
        rice[9][6] = 16'b00000_110000_11111;
        rice[9][7] = 16'b00000_110000_11111;
        rice[9][8] = 16'b00000_110000_11111;
        rice[9][9] = 16'b00000_110000_11111;
        rice[9][10] = 16'b00000_110000_11111;
        rice[9][11] = 16'b00000_110000_11111;
        rice[9][12] = 16'b00000_110000_11111;
        rice[9][13] = 16'b00000_000000_00000;
        rice[9][14] = 16'b00000_110000_11111;
        rice[10][0] = 16'b00000_110000_11111;
        rice[10][1] = 16'b00000_000000_00000;
        rice[10][2] = 16'b00000_000000_00000;
        rice[10][3] = 16'b00000_110000_11111;
        rice[10][4] = 16'b00000_110000_11111;
        rice[10][5] = 16'b00000_110000_11111;
        rice[10][6] = 16'b00000_110000_11111;
        rice[10][7] = 16'b00000_110000_11111;
        rice[10][8] = 16'b00000_110000_11111;
        rice[10][9] = 16'b00000_110000_11111;
        rice[10][10] = 16'b00000_110000_11111;
        rice[10][11] = 16'b00000_110000_11111;
        rice[10][12] = 16'b00000_000000_00000;
        rice[10][13] = 16'b00000_000000_00000;
        rice[10][14] = 16'b00000_110000_11111;
        rice[11][0] = 16'b00000_110000_11111;
        rice[11][1] = 16'b00000_000000_00000;
        rice[11][2] = 16'b00000_000000_00000;
        rice[11][3] = 16'b00000_110000_11111;
        rice[11][4] = 16'b00000_110000_11111;
        rice[11][5] = 16'b00000_110000_11111;
        rice[11][6] = 16'b00000_110000_11111;
        rice[11][7] = 16'b00000_110000_11111;
        rice[11][8] = 16'b00000_110000_11111;
        rice[11][9] = 16'b00000_110000_11111;
        rice[11][10] = 16'b00000_110000_11111;
        rice[11][11] = 16'b00000_110000_11111;
        rice[11][12] = 16'b00000_000000_00000;
        rice[11][13] = 16'b00000_000000_00000;
        rice[11][14] = 16'b00000_110000_11111;
        rice[12][0] = 16'b00000_110000_11111;
        rice[12][1] = 16'b00000_000000_00000;
        rice[12][2] = 16'b00000_000000_00000;
        rice[12][3] = 16'b00000_000000_00000;
        rice[12][4] = 16'b00000_000000_00000;
        rice[12][5] = 16'b00000_000000_00000;
        rice[12][6] = 16'b00000_110000_11111;
        rice[12][7] = 16'b00000_110000_11111;
        rice[12][8] = 16'b00000_110000_11111;
        rice[12][9] = 16'b00000_000000_00000;
        rice[12][10] = 16'b00000_000000_00000;
        rice[12][11] = 16'b00000_000000_00000;
        rice[12][12] = 16'b00000_000000_00000;
        rice[12][13] = 16'b00000_000000_00000;
        rice[12][14] = 16'b00000_110000_11111;
        rice[13][0] = 16'b00000_110000_11111;
        rice[13][1] = 16'b00000_000000_00000;
        rice[13][2] = 16'b00000_000000_00000;
        rice[13][3] = 16'b00000_000000_00000;
        rice[13][4] = 16'b00000_000000_00000;
        rice[13][5] = 16'b00000_000000_00000;
        rice[13][6] = 16'b00000_000000_00000;
        rice[13][7] = 16'b00000_000000_00000;
        rice[13][8] = 16'b00000_000000_00000;
        rice[13][9] = 16'b00000_000000_00000;
        rice[13][10] = 16'b00000_000000_00000;
        rice[13][11] = 16'b00000_000000_00000;
        rice[13][12] = 16'b00000_000000_00000;
        rice[13][13] = 16'b00000_000000_00000;
        rice[13][14] = 16'b00000_110000_11111;
        rice[14][0] = 16'b00000_110000_11111;
        rice[14][1] = 16'b00000_110000_11111;
        rice[14][2] = 16'b00000_110000_11111;
        rice[14][3] = 16'b00000_110000_11111;
        rice[14][4] = 16'b00000_110000_11111;
        rice[14][5] = 16'b00000_110000_11111;
        rice[14][6] = 16'b00000_110000_11111;
        rice[14][7] = 16'b00000_110000_11111;
        rice[14][8] = 16'b00000_110000_11111;
        rice[14][9] = 16'b00000_110000_11111;
        rice[14][10] = 16'b00000_110000_11111;
        rice[14][11] = 16'b00000_110000_11111;
        rice[14][12] = 16'b00000_110000_11111;
        rice[14][13] = 16'b00000_110000_11111;
        rice[14][14] = 16'b00000_110000_11111;
    
        
        tomato[0][0] = 16'b11001_000000_00000;
        tomato[0][1] = 16'b11001_000000_00000;
        tomato[0][2] = 16'b11001_000000_00000;
        tomato[0][3] = 16'b11001_000000_00000;
        tomato[0][4] = 16'b11001_000000_00000;
        tomato[0][5] = 16'b11001_000000_00000;
        tomato[0][6] = 16'b11001_000000_00000;
        tomato[0][7] = 16'b11001_000000_00000;
        tomato[0][8] = 16'b11001_000000_00000;
        tomato[0][9] = 16'b11001_000000_00000;
        tomato[0][10] = 16'b11001_000000_00000;
        tomato[0][11] = 16'b11001_000000_00000;
        tomato[0][12] = 16'b11001_000000_00000;
        tomato[0][13] = 16'b11001_000000_00000;
        tomato[0][14] = 16'b11001_000000_00000;
        tomato[1][0] = 16'b11001_000000_00000;
        tomato[1][1] = 16'b00000_000000_00000;
        tomato[1][2] = 16'b00000_000000_00000;
        tomato[1][3] = 16'b00000_000000_00000;
        tomato[1][4] = 16'b00000_000000_00000;
        tomato[1][5] = 16'b00000_000000_00000;
        tomato[1][6] = 16'b00000_000000_00000;
        tomato[1][7] = 16'b00000_000000_00000;
        tomato[1][8] = 16'b00000_000000_00000;
        tomato[1][9] = 16'b00000_000000_00000;
        tomato[1][10] = 16'b00000_000000_00000;
        tomato[1][11] = 16'b00000_000000_00000;
        tomato[1][12] = 16'b00000_000000_00000;
        tomato[1][13] = 16'b00000_000000_00000;
        tomato[1][14] = 16'b11001_000000_00000;
        tomato[2][0] = 16'b11001_000000_00000;
        tomato[2][1] = 16'b00000_000000_00000;
        tomato[2][2] = 16'b00000_000000_00000;
        tomato[2][3] = 16'b00000_000000_00000;
        tomato[2][4] = 16'b00000_011100_00000;
        tomato[2][5] = 16'b00000_011100_00000;
        tomato[2][6] = 16'b00000_011100_00000;
        tomato[2][7] = 16'b11001_000000_00000;
        tomato[2][8] = 16'b00000_011100_00000;
        tomato[2][9] = 16'b00000_011100_00000;
        tomato[2][10] = 16'b00000_011100_00000;
        tomato[2][11] = 16'b00000_000000_00000;
        tomato[2][12] = 16'b00000_000000_00000;
        tomato[2][13] = 16'b00000_000000_00000;
        tomato[2][14] = 16'b11001_000000_00000;
        tomato[3][0] = 16'b11001_000000_00000;
        tomato[3][1] = 16'b00000_000000_00000;
        tomato[3][2] = 16'b00000_000000_00000;
        tomato[3][3] = 16'b00000_000000_00000;
        tomato[3][4] = 16'b11001_000000_00000;
        tomato[3][5] = 16'b11001_000000_00000;
        tomato[3][6] = 16'b00000_011100_00000;
        tomato[3][7] = 16'b00000_011100_00000;
        tomato[3][8] = 16'b00000_011100_00000;
        tomato[3][9] = 16'b11001_000000_00000;
        tomato[3][10] = 16'b11001_000000_00000;
        tomato[3][11] = 16'b00000_000000_00000;
        tomato[3][12] = 16'b00000_000000_00000;
        tomato[3][13] = 16'b00000_000000_00000;
        tomato[3][14] = 16'b11001_000000_00000;
        tomato[4][0] = 16'b11001_000000_00000;
        tomato[4][1] = 16'b00000_000000_00000;
        tomato[4][2] = 16'b00000_000000_00000;
        tomato[4][3] = 16'b11001_000000_00000;
        tomato[4][4] = 16'b00000_011100_00000;
        tomato[4][5] = 16'b00000_011100_00000;
        tomato[4][6] = 16'b11001_000000_00000;
        tomato[4][7] = 16'b11001_000000_00000;
        tomato[4][8] = 16'b11001_000000_00000;
        tomato[4][9] = 16'b00000_011100_00000;
        tomato[4][10] = 16'b00000_011100_00000;
        tomato[4][11] = 16'b11001_000000_00000;
        tomato[4][12] = 16'b00000_000000_00000;
        tomato[4][13] = 16'b00000_000000_00000;
        tomato[4][14] = 16'b11001_000000_00000;
        tomato[5][0] = 16'b11001_000000_00000;
        tomato[5][1] = 16'b00000_000000_00000;
        tomato[5][2] = 16'b11001_000000_00000;
        tomato[5][3] = 16'b00000_011100_00000;
        tomato[5][4] = 16'b00000_011100_00000;
        tomato[5][5] = 16'b11001_000000_00000;
        tomato[5][6] = 16'b11001_000000_00000;
        tomato[5][7] = 16'b11001_000000_00000;
        tomato[5][8] = 16'b11001_000000_00000;
        tomato[5][9] = 16'b11001_000000_00000;
        tomato[5][10] = 16'b00000_011100_00000;
        tomato[5][11] = 16'b00000_011100_00000;
        tomato[5][12] = 16'b11001_000000_00000;
        tomato[5][13] = 16'b00000_000000_00000;
        tomato[5][14] = 16'b11001_000000_00000;
        tomato[6][0] = 16'b11001_000000_00000;
        tomato[6][1] = 16'b00000_000000_00000;
        tomato[6][2] = 16'b11001_000000_00000;
        tomato[6][3] = 16'b11001_000000_00000;
        tomato[6][4] = 16'b11001_000000_00000;
        tomato[6][5] = 16'b11001_000000_00000;
        tomato[6][6] = 16'b11001_000000_00000;
        tomato[6][7] = 16'b11001_000000_00000;
        tomato[6][8] = 16'b11001_000000_00000;
        tomato[6][9] = 16'b11001_000000_00000;
        tomato[6][10] = 16'b11001_000000_00000;
        tomato[6][11] = 16'b11001_000000_00000;
        tomato[6][12] = 16'b11001_000000_00000;
        tomato[6][13] = 16'b00000_000000_00000;
        tomato[6][14] = 16'b11001_000000_00000;
        tomato[7][0] = 16'b11001_000000_00000;
        tomato[7][1] = 16'b00000_000000_00000;
        tomato[7][2] = 16'b11001_000000_00000;
        tomato[7][3] = 16'b11001_000000_00000;
        tomato[7][4] = 16'b11001_000000_00000;
        tomato[7][5] = 16'b11001_000000_00000;
        tomato[7][6] = 16'b11001_000000_00000;
        tomato[7][7] = 16'b11001_000000_00000;
        tomato[7][8] = 16'b11001_000000_00000;
        tomato[7][9] = 16'b11001_000000_00000;
        tomato[7][10] = 16'b11001_000000_00000;
        tomato[7][11] = 16'b11001_000000_00000;
        tomato[7][12] = 16'b11001_000000_00000;
        tomato[7][13] = 16'b00000_000000_00000;
        tomato[7][14] = 16'b11001_000000_00000;
        tomato[8][0] = 16'b11001_000000_00000;
        tomato[8][1] = 16'b00000_000000_00000;
        tomato[8][2] = 16'b11001_000000_00000;
        tomato[8][3] = 16'b11001_000000_00000;
        tomato[8][4] = 16'b11001_000000_00000;
        tomato[8][5] = 16'b11001_000000_00000;
        tomato[8][6] = 16'b11001_000000_00000;
        tomato[8][7] = 16'b11001_000000_00000;
        tomato[8][8] = 16'b11001_000000_00000;
        tomato[8][9] = 16'b11001_000000_00000;
        tomato[8][10] = 16'b11001_000000_00000;
        tomato[8][11] = 16'b11001_000000_00000;
        tomato[8][12] = 16'b11001_000000_00000;
        tomato[8][13] = 16'b00000_000000_00000;
        tomato[8][14] = 16'b11001_000000_00000;
        tomato[9][0] = 16'b11001_000000_00000;
        tomato[9][1] = 16'b00000_000000_00000;
        tomato[9][2] = 16'b11001_000000_00000;
        tomato[9][3] = 16'b11001_000000_00000;
        tomato[9][4] = 16'b11001_000000_00000;
        tomato[9][5] = 16'b11001_000000_00000;
        tomato[9][6] = 16'b11001_000000_00000;
        tomato[9][7] = 16'b11001_000000_00000;
        tomato[9][8] = 16'b11001_000000_00000;
        tomato[9][9] = 16'b11001_000000_00000;
        tomato[9][10] = 16'b11001_000000_00000;
        tomato[9][11] = 16'b11001_000000_00000;
        tomato[9][12] = 16'b11001_000000_00000;
        tomato[9][13] = 16'b00000_000000_00000;
        tomato[9][14] = 16'b11001_000000_00000;
        tomato[10][0] = 16'b11001_000000_00000;
        tomato[10][1] = 16'b00000_000000_00000;
        tomato[10][2] = 16'b10001_000000_00000;
        tomato[10][3] = 16'b11001_000000_00000;
        tomato[10][4] = 16'b11001_000000_00000;
        tomato[10][5] = 16'b11001_000000_00000;
        tomato[10][6] = 16'b11001_000000_00000;
        tomato[10][7] = 16'b11001_000000_00000;
        tomato[10][8] = 16'b11001_000000_00000;
        tomato[10][9] = 16'b11001_000000_00000;
        tomato[10][10] = 16'b11001_000000_00000;
        tomato[10][11] = 16'b11001_000000_00000;
        tomato[10][12] = 16'b10001_000000_00000;
        tomato[10][13] = 16'b00000_000000_00000;
        tomato[10][14] = 16'b11001_000000_00000;
        tomato[11][0] = 16'b11001_000000_00000;
        tomato[11][1] = 16'b00000_000000_00000;
        tomato[11][2] = 16'b00000_000000_00000;
        tomato[11][3] = 16'b10001_000000_00000;
        tomato[11][4] = 16'b10001_000000_00000;
        tomato[11][5] = 16'b10001_000000_00000;
        tomato[11][6] = 16'b11001_000000_00000;
        tomato[11][7] = 16'b11001_000000_00000;
        tomato[11][8] = 16'b11001_000000_00000;
        tomato[11][9] = 16'b10001_000000_00000;
        tomato[11][10] = 16'b10001_000000_00000;
        tomato[11][11] = 16'b10001_000000_00000;
        tomato[11][12] = 16'b00000_000000_00000;
        tomato[11][13] = 16'b00000_000000_00000;
        tomato[11][14] = 16'b11001_000000_00000;
        tomato[12][0] = 16'b11001_000000_00000;
        tomato[12][1] = 16'b00000_000000_00000;
        tomato[12][2] = 16'b00000_000000_00000;
        tomato[12][3] = 16'b00000_000000_00000;
        tomato[12][4] = 16'b00000_000000_00000;
        tomato[12][5] = 16'b10001_000000_00000;
        tomato[12][6] = 16'b10001_000000_00000;
        tomato[12][7] = 16'b10001_000000_00000;
        tomato[12][8] = 16'b10001_000000_00000;
        tomato[12][9] = 16'b10001_000000_00000;
        tomato[12][10] = 16'b00000_000000_00000;
        tomato[12][11] = 16'b00000_000000_00000;
        tomato[12][12] = 16'b00000_000000_00000;
        tomato[12][13] = 16'b00000_000000_00000;
        tomato[12][14] = 16'b11001_000000_00000;
        tomato[13][0] = 16'b11001_000000_00000;
        tomato[13][1] = 16'b00000_000000_00000;
        tomato[13][2] = 16'b00000_000000_00000;
        tomato[13][3] = 16'b00000_000000_00000;
        tomato[13][4] = 16'b00000_000000_00000;
        tomato[13][5] = 16'b00000_000000_00000;
        tomato[13][6] = 16'b00000_000000_00000;
        tomato[13][7] = 16'b00000_000000_00000;
        tomato[13][8] = 16'b00000_000000_00000;
        tomato[13][9] = 16'b00000_000000_00000;
        tomato[13][10] = 16'b00000_000000_00000;
        tomato[13][11] = 16'b00000_000000_00000;
        tomato[13][12] = 16'b00000_000000_00000;
        tomato[13][13] = 16'b00000_000000_00000;
        tomato[13][14] = 16'b11001_000000_00000;
        tomato[14][0] = 16'b11001_000000_00000;
        tomato[14][1] = 16'b11001_000000_00000;
        tomato[14][2] = 16'b11001_000000_00000;
        tomato[14][3] = 16'b11001_000000_00000;
        tomato[14][4] = 16'b11001_000000_00000;
        tomato[14][5] = 16'b11001_000000_00000;
        tomato[14][6] = 16'b11001_000000_00000;
        tomato[14][7] = 16'b11001_000000_00000;
        tomato[14][8] = 16'b11001_000000_00000;
        tomato[14][9] = 16'b11001_000000_00000;
        tomato[14][10] = 16'b11001_000000_00000;
        tomato[14][11] = 16'b11001_000000_00000;
        tomato[14][12] = 16'b11001_000000_00000;
        tomato[14][13] = 16'b11001_000000_00000;
        tomato[14][14] = 16'b11001_000000_00000;
        
        chicken[0][0] = 16'b11111_101111_01111;
        chicken[0][1] = 16'b11111_101111_01111;
        chicken[0][2] = 16'b11111_101111_01111;
        chicken[0][3] = 16'b11111_101111_01111;
        chicken[0][4] = 16'b11111_101111_01111;
        chicken[0][5] = 16'b11111_101111_01111;
        chicken[0][6] = 16'b11111_101111_01111;
        chicken[0][7] = 16'b11111_101111_01111;
        chicken[0][8] = 16'b11111_101111_01111;
        chicken[0][9] = 16'b11111_101111_01111;
        chicken[0][10] = 16'b11111_101111_01111;
        chicken[0][11] = 16'b11111_101111_01111;
        chicken[0][12] = 16'b11111_101111_01111;
        chicken[0][13] = 16'b11111_101111_01111;
        chicken[0][14] = 16'b11111_101111_01111;
        chicken[1][0] = 16'b11111_101111_01111;
        chicken[1][1] = 16'b00000_000000_00000;
        chicken[1][2] = 16'b00000_000000_00000;
        chicken[1][3] = 16'b00000_000000_00000;
        chicken[1][4] = 16'b00000_000000_00000;
        chicken[1][5] = 16'b00000_000000_00000;
        chicken[1][6] = 16'b00000_000000_00000;
        chicken[1][7] = 16'b00000_000000_00000;
        chicken[1][8] = 16'b00000_000000_00000;
        chicken[1][9] = 16'b11111_101000_00100;
        chicken[1][10] = 16'b11111_101000_00100;
        chicken[1][11] = 16'b11111_101000_00100;
        chicken[1][12] = 16'b00000_000000_00000;
        chicken[1][13] = 16'b00000_000000_00000;
        chicken[1][14] = 16'b11111_101111_01111;
        chicken[2][0] = 16'b11111_101111_01111;
        chicken[2][1] = 16'b00000_000000_00000;
        chicken[2][2] = 16'b00000_000000_00000;
        chicken[2][3] = 16'b00000_000000_00000;
        chicken[2][4] = 16'b00000_000000_00000;
        chicken[2][5] = 16'b00000_000000_00000;
        chicken[2][6] = 16'b00000_000000_00000;
        chicken[2][7] = 16'b11111_101000_00100;
        chicken[2][8] = 16'b11111_101000_00100;
        chicken[2][9] = 16'b11111_101111_01111;
        chicken[2][10] = 16'b11111_101111_01111;
        chicken[2][11] = 16'b11111_101111_01111;
        chicken[2][12] = 16'b11111_101000_00100;
        chicken[2][13] = 16'b00000_000000_00000;
        chicken[2][14] = 16'b11111_101111_01111;
        chicken[3][0] = 16'b11111_101111_01111;
        chicken[3][1] = 16'b00000_000000_00000;
        chicken[3][2] = 16'b00000_000000_00000;
        chicken[3][3] = 16'b00000_000000_00000;
        chicken[3][4] = 16'b00000_000000_00000;
        chicken[3][5] = 16'b00000_000000_00000;
        chicken[3][6] = 16'b00000_000000_00000;
        chicken[3][7] = 16'b11111_101000_00100;
        chicken[3][8] = 16'b11111_101111_01111;
        chicken[3][9] = 16'b11111_101111_01111;
        chicken[3][10] = 16'b11111_101111_01111;
        chicken[3][11] = 16'b11111_101111_01111;
        chicken[3][12] = 16'b11111_101000_00100;
        chicken[3][13] = 16'b11111_101000_00100;
        chicken[3][14] = 16'b11111_101111_01111;
        chicken[4][0] = 16'b11111_101111_01111;
        chicken[4][1] = 16'b00000_000000_00000;
        chicken[4][2] = 16'b00000_000000_00000;
        chicken[4][3] = 16'b00000_000000_00000;
        chicken[4][4] = 16'b00000_000000_00000;
        chicken[4][5] = 16'b00000_000000_00000;
        chicken[4][6] = 16'b11111_101000_00100;
        chicken[4][7] = 16'b11111_101111_01111;
        chicken[4][8] = 16'b11111_101111_01111;
        chicken[4][9] = 16'b11111_101111_01111;
        chicken[4][10] = 16'b11111_101111_01111;
        chicken[4][11] = 16'b11111_101111_01111;
        chicken[4][12] = 16'b11111_101111_01111;
        chicken[4][13] = 16'b11111_101000_00100;
        chicken[4][14] = 16'b11111_101111_01111;
        chicken[5][0] = 16'b11111_101111_01111;
        chicken[5][1] = 16'b00000_000000_00000;
        chicken[5][2] = 16'b00000_000000_00000;
        chicken[5][3] = 16'b00000_000000_00000;
        chicken[5][4] = 16'b00000_000000_00000;
        chicken[5][5] = 16'b00000_000000_00000;
        chicken[5][6] = 16'b11111_101000_00100;
        chicken[5][7] = 16'b11111_101111_01111;
        chicken[5][8] = 16'b11111_101111_01111;
        chicken[5][9] = 16'b11111_101111_01111;
        chicken[5][10] = 16'b11111_101111_01111;
        chicken[5][11] = 16'b11111_101111_01111;
        chicken[5][12] = 16'b11111_101000_00100;
        chicken[5][13] = 16'b11111_101000_00100;
        chicken[5][14] = 16'b11111_101111_01111;
        chicken[6][0] = 16'b11111_101111_01111;
        chicken[6][1] = 16'b00000_000000_00000;
        chicken[6][2] = 16'b00000_000000_00000;
        chicken[6][3] = 16'b00000_000000_00000;
        chicken[6][4] = 16'b00000_000000_00000;
        chicken[6][5] = 16'b00000_000000_00000;
        chicken[6][6] = 16'b11111_101000_00100;
        chicken[6][7] = 16'b11111_101111_01111;
        chicken[6][8] = 16'b11111_101111_01111;
        chicken[6][9] = 16'b11111_101111_01111;
        chicken[6][10] = 16'b11111_101111_01111;
        chicken[6][11] = 16'b11111_101111_01111;
        chicken[6][12] = 16'b11111_101000_00100;
        chicken[6][13] = 16'b00000_000000_00000;
        chicken[6][14] = 16'b11111_101111_01111;
        chicken[7][0] = 16'b11111_101111_01111;
        chicken[7][1] = 16'b00000_000000_00000;
        chicken[7][2] = 16'b00000_000000_00000;
        chicken[7][3] = 16'b00000_000000_00000;
        chicken[7][4] = 16'b00000_000000_00000;
        chicken[7][5] = 16'b11111_101000_00100;
        chicken[7][6] = 16'b11111_101111_01111;
        chicken[7][7] = 16'b11111_101111_01111;
        chicken[7][8] = 16'b11111_101111_01111;
        chicken[7][9] = 16'b11111_101111_01111;
        chicken[7][10] = 16'b11111_101111_01111;
        chicken[7][11] = 16'b11111_101000_00100;
        chicken[7][12] = 16'b11111_101000_00100;
        chicken[7][13] = 16'b00000_000000_00000;
        chicken[7][14] = 16'b11111_101111_01111;
        chicken[8][0] = 16'b11111_101111_01111;
        chicken[8][1] = 16'b00000_000000_00000;
        chicken[8][2] = 16'b00000_000000_00000;
        chicken[8][3] = 16'b00000_000000_00000;
        chicken[8][4] = 16'b00000_000000_00000;
        chicken[8][5] = 16'b11111_101000_00100;
        chicken[8][6] = 16'b11111_101111_01111;
        chicken[8][7] = 16'b11111_101111_01111;
        chicken[8][8] = 16'b11111_101111_01111;
        chicken[8][9] = 16'b11111_101000_00100;
        chicken[8][10] = 16'b11111_101000_00100;
        chicken[8][11] = 16'b11111_101000_00100;
        chicken[8][12] = 16'b00000_000000_00000;
        chicken[8][13] = 16'b00000_000000_00000;
        chicken[8][14] = 16'b11111_101111_01111;
        chicken[9][0] = 16'b11111_101111_01111;
        chicken[9][1] = 16'b00000_000000_00000;
        chicken[9][2] = 16'b00000_000000_00000;
        chicken[9][3] = 16'b00000_000000_00000;
        chicken[9][4] = 16'b11111_101000_00100;
        chicken[9][5] = 16'b11111_101111_01111;
        chicken[9][6] = 16'b11111_101111_01111;
        chicken[9][7] = 16'b11111_101000_00100;
        chicken[9][8] = 16'b11111_101000_00100;
        chicken[9][9] = 16'b00000_000000_00000;
        chicken[9][10] = 16'b00000_000000_00000;
        chicken[9][11] = 16'b00000_000000_00000;
        chicken[9][12] = 16'b00000_000000_00000;
        chicken[9][13] = 16'b00000_000000_00000;
        chicken[9][14] = 16'b11111_101111_01111;
        chicken[10][0] = 16'b11111_101111_01111;
        chicken[10][1] = 16'b00000_000000_00000;
        chicken[10][2] = 16'b00000_000000_00000;
        chicken[10][3] = 16'b11111_111110_11111;
        chicken[10][4] = 16'b11111_101000_00100;
        chicken[10][5] = 16'b11111_101000_00100;
        chicken[10][6] = 16'b11111_101000_00100;
        chicken[10][7] = 16'b00000_000000_00000;
        chicken[10][8] = 16'b00000_000000_00000;
        chicken[10][9] = 16'b00000_000000_00000;
        chicken[10][10] = 16'b00000_000000_00000;
        chicken[10][11] = 16'b00000_000000_00000;
        chicken[10][12] = 16'b00000_000000_00000;
        chicken[10][13] = 16'b00000_000000_00000;
        chicken[10][14] = 16'b11111_101111_01111;
        chicken[11][0] = 16'b11111_101111_01111;
        chicken[11][1] = 16'b00000_000000_00000;
        chicken[11][2] = 16'b11111_111110_11111;
        chicken[11][3] = 16'b11111_111110_11111;
        chicken[11][4] = 16'b11111_111110_11111;
        chicken[11][5] = 16'b00000_000000_00000;
        chicken[11][6] = 16'b00000_000000_00000;
        chicken[11][7] = 16'b00000_000000_00000;
        chicken[11][8] = 16'b00000_000000_00000;
        chicken[11][9] = 16'b00000_000000_00000;
        chicken[11][10] = 16'b00000_000000_00000;
        chicken[11][11] = 16'b00000_000000_00000;
        chicken[11][12] = 16'b00000_000000_00000;
        chicken[11][13] = 16'b00000_000000_00000;
        chicken[11][14] = 16'b11111_101111_01111;
        chicken[12][0] = 16'b11111_101111_01111;
        chicken[12][1] = 16'b11111_111110_11111;
        chicken[12][2] = 16'b11111_111110_11111;
        chicken[12][3] = 16'b11111_111110_11111;
        chicken[12][4] = 16'b00000_000000_00000;
        chicken[12][5] = 16'b00000_000000_00000;
        chicken[12][6] = 16'b00000_000000_00000;
        chicken[12][7] = 16'b00000_000000_00000;
        chicken[12][8] = 16'b00000_000000_00000;
        chicken[12][9] = 16'b00000_000000_00000;
        chicken[12][10] = 16'b00000_000000_00000;
        chicken[12][11] = 16'b00000_000000_00000;
        chicken[12][12] = 16'b00000_000000_00000;
        chicken[12][13] = 16'b00000_000000_00000;
        chicken[12][14] = 16'b11111_101111_01111;
        chicken[13][0] = 16'b11111_101111_01111;
        chicken[13][1] = 16'b11111_111110_11111;
        chicken[13][2] = 16'b11111_111110_11111;
        chicken[13][3] = 16'b00000_000000_00000;
        chicken[13][4] = 16'b00000_000000_00000;
        chicken[13][5] = 16'b00000_000000_00000;
        chicken[13][6] = 16'b00000_000000_00000;
        chicken[13][7] = 16'b00000_000000_00000;
        chicken[13][8] = 16'b00000_000000_00000;
        chicken[13][9] = 16'b00000_000000_00000;
        chicken[13][10] = 16'b00000_000000_00000;
        chicken[13][11] = 16'b00000_000000_00000;
        chicken[13][12] = 16'b00000_000000_00000;
        chicken[13][13] = 16'b00000_000000_00000;
        chicken[13][14] = 16'b11111_101111_01111;
        chicken[14][0] = 16'b11111_101111_01111;
        chicken[14][1] = 16'b11111_101111_01111;
        chicken[14][2] = 16'b11111_101111_01111;
        chicken[14][3] = 16'b11111_101111_01111;
        chicken[14][4] = 16'b11111_101111_01111;
        chicken[14][5] = 16'b11111_101111_01111;
        chicken[14][6] = 16'b11111_101111_01111;
        chicken[14][7] = 16'b11111_101111_01111;
        chicken[14][8] = 16'b11111_101111_01111;
        chicken[14][9] = 16'b11111_101111_01111;
        chicken[14][10] = 16'b11111_101111_01111;
        chicken[14][11] = 16'b11111_101111_01111;
        chicken[14][12] = 16'b11111_101111_01111;
        chicken[14][13] = 16'b11111_101111_01111;
        chicken[14][14] = 16'b11111_101111_01111;

        
    end
    
    always @(posedge clk_25MHz) begin
        if (x >= ONION_TOP_LEFT_X && x < ONION_TOP_LEFT_X+15 && y >= ONION_TOP_LEFT_Y && y < ONION_TOP_LEFT_Y+15) begin
            oled_data <= onion[y - ONION_TOP_LEFT_Y][x - ONION_TOP_LEFT_X]; // offset your image to screen position
        end 
        else if (x >= RICE_TOP_LEFT_X && x < RICE_TOP_LEFT_X+15 && y >= RICE_TOP_LEFT_Y && y < RICE_TOP_LEFT_Y+15) begin
            oled_data <= rice[y - RICE_TOP_LEFT_Y][x - RICE_TOP_LEFT_X]; // offset your image to screen position
        end         
        else if (x >= CHICKEN_TOP_LEFT_X && x < CHICKEN_TOP_LEFT_X+15 && y >= CHICKEN_TOP_LEFT_Y && y < CHICKEN_TOP_LEFT_Y+15) begin
            oled_data <= chicken[y - CHICKEN_TOP_LEFT_Y][x - CHICKEN_TOP_LEFT_X]; // offset your image to screen position
        end         
        else if (x >= TOMATO_TOP_LEFT_X && x < TOMATO_TOP_LEFT_X+15 && y >= TOMATO_TOP_LEFT_Y && y < TOMATO_TOP_LEFT_Y+15) begin
            oled_data <= tomato[y - TOMATO_TOP_LEFT_Y][x - TOMATO_TOP_LEFT_X]; // offset your image to screen position
        end 
        else begin
            oled_data <= 0;
        end
    end

endmodule
